--Copyright (C)2014-2025 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.11.01 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Thu May 15 12:11:11 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_basic is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_basic;

architecture Behavioral of Gowin_pROM_basic is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C6992B653CAFBD8E603210F816852222834CC0D81110D2134F3554400C1B1282",
            INIT_RAM_01 => X"C64939556CEAE29F59569B269A244222266662262260AF12422B9C125F34D509",
            INIT_RAM_02 => X"CAEBAD29B2AAD1C889F6944B26C2598C21E85714F9C1E8E9692B548A459F57B2",
            INIT_RAM_03 => X"4E4F704B96008829697A7C896DCC6EEAA9BABEB553DD5B356B32D5A568AE5AEE",
            INIT_RAM_04 => X"6259D1CF297E8995124709D1894A4A55696C81D3D259BFFFADDD081C931D3FFF",
            INIT_RAM_05 => X"E354D453A65A765AA553295F5347348F593A2D91D4A6F278B4E7344DE6629346",
            INIT_RAM_06 => X"812C006403626D13128020451B2EA4200567420235C716B954ACD4666311BE2C",
            INIT_RAM_07 => X"402FE67406919878DEB782525C9A40128214A4F175F7935F50AC32D0440A6C52",
            INIT_RAM_08 => X"4E0EA95529839D1E517918381EBB4BB4B478850DE069918B2100200093D3F39C",
            INIT_RAM_09 => X"5835722CD2019949488EF39128654D239331924B22E25C006A0C860050776A89",
            INIT_RAM_0A => X"1DFC04A00251B8CCE64CD2091852BADECC084055053A891C6F910A4933244198",
            INIT_RAM_0B => X"08A5210504A499050025080C02A0828849ABA0A50FC472AA11908801A1000828",
            INIT_RAM_0C => X"4E380331422168861ACD1E966B08440990A44A75049998DC8686A940CC01E29A",
            INIT_RAM_0D => X"A4435DA80A64721001E4FDBCE965013895FE46232D7609CE5395A8ED30CDA800",
            INIT_RAM_0E => X"C90DC690B110A82204004F6800311949A0A1D8F5406DFCA00109095DA2D2B056",
            INIT_RAM_0F => X"48344D040428C83A2410200800C223A9AEA728264C1A39805C80C124D0230041",
            INIT_RAM_10 => X"F493151694931246687B66C0301004824A1617A81E2430D0CE8A051543989CAC",
            INIT_RAM_11 => X"8107324E8A449A76736552282C551D0C694A7FC68B49000F4B0C03AE74258944",
            INIT_RAM_12 => X"8C046D0218E71237912234A540A2AD1EBB0A8E51649A09448853FE186958AE45",
            INIT_RAM_13 => X"B25A641965834E12B784E9DD0444A46189E5985977EEECB40008250952479CEF",
            INIT_RAM_14 => X"8E4820808861C5205B295094A5225C1A45A1AF103224E64C6C91DAA696C7AB2C",
            INIT_RAM_15 => X"42530DA4458102D68A08A24666A5301C452F0BCD84140B410388062814740010",
            INIT_RAM_16 => X"A508BD46CF12494910A8B101025888A4E61109E33204C62D406BB65FADF09FF4",
            INIT_RAM_17 => X"12A17010782800090C264D225693339BB9350041445504C6EE1E09541D561860",
            INIT_RAM_18 => X"AC821667590CA7EAEA164C832E9011E7449004A3D8D0B8CEBC215AE3E3414080",
            INIT_RAM_19 => X"2434B4280E521DD074E7A8A5427849D90CB3260363834BE0CB0EA14C8128C82A",
            INIT_RAM_1A => X"63C65916B4855C8CB24AC940426148930015E82D53122000DD1433B41015CD58",
            INIT_RAM_1B => X"048205A02C0A103EBAA005023D244C0A4C83119C488222221652CA32E7994462",
            INIT_RAM_1C => X"08501301A272411330F4C080000020F080952C8E24266407930480000480C095",
            INIT_RAM_1D => X"2D938F18A2930891922244A822B281451006212C03C830AEF11C052235E34724",
            INIT_RAM_1E => X"E977A5745549581038418702B187AEADC12452060100FBB19AA10028711164C4",
            INIT_RAM_1F => X"7661008A88483050412810103BFBBFBAE88823FB044715FD5FD4E8A41410069D",
            INIT_RAM_20 => X"2BAAD2B490110AFEAFE8B402B4AD3BAE56C1002D03002AC48303AF901405A908",
            INIT_RAM_21 => X"C2BFABF80221868A00A032B7916CA2D200A5020A62D3EB4235BC15D4304304BD",
            INIT_RAM_22 => X"A568504911675A6A199B868B114022CA1CBA729C804101C2B1C31C246F5F5200",
            INIT_RAM_23 => X"9112E251A1CD5920223133918CAC8E901BB3F4898711450C733A118118DAE946",
            INIT_RAM_24 => X"B0990CD094B3976058A001007E06065297830404C8B13998A520880CA2D51204",
            INIT_RAM_25 => X"506B15A070763F07432504026ACAD76497F9206913800EA649E506E000D7FB5F",
            INIT_RAM_26 => X"42106B18302F060D0D1B351A4B2EE6B724E11281089C616F01E4E98002052032",
            INIT_RAM_27 => X"252B02649D3504D5CBCA2102062CA2880851AE7D55B5D4D8D8483573FD7B6010",
            INIT_RAM_28 => X"94D01298251582509419524051484A424142CE86610C082C822255E3F10E0406",
            INIT_RAM_29 => X"86030321800248493C10C079E90082C208888044488524B1123C76425A50B086",
            INIT_RAM_2A => X"884E74821547812A46A014EC88815B140D012144AD0D1B4A96330724884397A4",
            INIT_RAM_2B => X"549C9A990A520722108E440B598466863840D61E3071F4A01B29136D44EEFED9",
            INIT_RAM_2C => X"BD2980CA0E1253016208704EC0115E32B05204D26484869ED94B231526A45396",
            INIT_RAM_2D => X"B4A5749A604E14645108C80A078A821457DCA5B4BE235F5DA7100FA286BE4B21",
            INIT_RAM_2E => X"2126E3056240C0216A41B0142BC8EC9A942A52624116B50580088D290785D992",
            INIT_RAM_2F => X"05DC202D898AD18EDA16804256903520A91002140A55B1252A216A1E46260332",
            INIT_RAM_30 => X"544012FE2810308921062085C80838905090800818B2890E0104289301CECA05",
            INIT_RAM_31 => X"B0206B20A06A80205C0C11D0E08A682006982C02872AFD290428CB09A2024978",
            INIT_RAM_32 => X"06D2444000009400901040C7044A68A0C002A8483100543076190E4EC310C104",
            INIT_RAM_33 => X"C39900669661CF037494A5AA3B643B4B9B9BB00B202278D9109A03024A407514",
            INIT_RAM_34 => X"2000E12A20910909948820A9BCD87A20F14D4249042124103C3482006032E821",
            INIT_RAM_35 => X"8BC534904248A6B1192103925925B5622B1722859723000151D0016CEC8C6700",
            INIT_RAM_36 => X"4294624283E81043A0CC1143F4218C912890E48681AE2DFB79C00A12D2731274",
            INIT_RAM_37 => X"6FC025CD5D84060D10224244E29088271AAA233200303C222C75000D4C0B0130",
            INIT_RAM_38 => X"788D26246D88EBCA8087E4BB46A5C5B112093041326048706D801E81F008FC40",
            INIT_RAM_39 => X"301094A8026220816AD272566C2304368E418490939135BDA12C24190910AFED",
            INIT_RAM_3A => X"46636A500264C2262A656B138CA80150140141080000806254144E0820405792",
            INIT_RAM_3B => X"C09ED2444C04936E142A0244294284130307405183021C0CB6481810B2204202",
            INIT_RAM_3C => X"61309413023A6A1502E2310188610221449781282100090809B7C9443C12D281",
            INIT_RAM_3D => X"36DD14BCD309672F108318822A4473493496F20D14A12B6218C8D51001002A2A",
            INIT_RAM_3E => X"4D1A442480B4409B294094B0988825B5400C8B12D90114310941AD34D14BD84A",
            INIT_RAM_3F => X"D11644AB62CB0F0D13413B30CFD1FC08860B6496C49689DEA9DA104440A0281B"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"34590643AA699C8B65A110116970D31D7D92732E7BB52EE5A00000E125929190",
            INIT_RAM_01 => X"8EAA9A2AA43A9C6ED6B6040A201E8511515151551540C600114D18DAC0B2FBF8",
            INIT_RAM_02 => X"A0C335CA21C21AFDC42A59822B1BF80A45C5644978CEE7B2E75D170BC94B669A",
            INIT_RAM_03 => X"0BBA89048B052F215EFD776EA19BA38022D6634A01A29A34F0114D4068077EC6",
            INIT_RAM_04 => X"21A4A08085B04098846A8CA2CC326190C48D8E68B7A2F5D0A8E3DD396575CA2A",
            INIT_RAM_05 => X"992B9A644E68360700F3354402821A5A86211E8A04C9863B610200C6E22C45E2",
            INIT_RAM_06 => X"93CD01400A2648705BC40440060007624A1B4190400E0930D988A42265998534",
            INIT_RAM_07 => X"58C1422C0414435084240000154200C5C01D1424A80500220525A04146BF0432",
            INIT_RAM_08 => X"E000108752092A421702C745808AA8882A0800244502A57246202080A2D90141",
            INIT_RAM_09 => X"1020A128A10150790088A25068A1108A882A024800A411020C5854020A802082",
            INIT_RAM_0A => X"08A882038D154E0A020890081A2404B48041020025000830CA21D46151404542",
            INIT_RAM_0B => X"028501D400A4006C24890ED52A0900C00AAAB0254AA940A258C2084004484103",
            INIT_RAM_0C => X"C9DA3484106D4894400812A003540448142492646145511510948B098B094400",
            INIT_RAM_0D => X"800050085220D81ACD4204200C4C904200888C262200C000210008508D0B6A76",
            INIT_RAM_0E => X"080C4E540464150829448000A43502544C9885083F02291548C9044400108450",
            INIT_RAM_0F => X"083640160752B2222055010004015509514828A80112208001008582008A0005",
            INIT_RAM_10 => X"96D016084ED01251465A02908204549008A190084444251208E025144A8915A8",
            INIT_RAM_11 => X"599110961160102AA23002342A51CD5C0400D5310C04A4292AA0558923252A6C",
            INIT_RAM_12 => X"00410246820830A13608888068A0788EA80A4814201000924006A914C24E9EC9",
            INIT_RAM_13 => X"055A24824042101C31000945B7B1A66916B454310012A000051DBCB140402008",
            INIT_RAM_14 => X"8252A8882108088000909036A0000442344D08510A00A88A9AA050B690615009",
            INIT_RAM_15 => X"421B004900081024C220225141822C04144A12BB08451345209D1088A0010414",
            INIT_RAM_16 => X"A06A4202028B4B616A2C0420689566E000174A9004505890D8155615088508A1",
            INIT_RAM_17 => X"80FA88040000020E2290080004A82200A881040544040A808214088000141380",
            INIT_RAM_18 => X"2008233281442010052001004614000B440400023081228520BA940502020000",
            INIT_RAM_19 => X"9D090401400120802154136019084441D3AA0801C27A921849440147B7018010",
            INIT_RAM_1A => X"06149825B54046082052D016C697640119A040A1204AD9710001202387A831A4",
            INIT_RAM_1B => X"04008130018C0251064B0718480A084A89F20185A11444440410922004108000",
            INIT_RAM_1C => X"0EA041120001421050A880B04001B6A081A1495420A834701004B12846888205",
            INIT_RAM_1D => X"000180A800130E4180210E4F9390454420121544800200A220005C8080420014",
            INIT_RAM_1E => X"522400A10544400C151000EC913155220620A8680EDFAA8A88500080102A0000",
            INIT_RAM_1F => X"73E005F56404011440EDDCCC90411555515F98285EA9AAA800090002AEFD86A0",
            INIT_RAM_20 => X"4554A108A52BF554000075142000014252430C0900441A0422440815180421BA",
            INIT_RAM_21 => X"05550002AF58102002A2845008253426409DB43360A56800040022A820000502",
            INIT_RAM_22 => X"080282007A1034C505609698243848342154A420B921904451410428600AA1FC",
            INIT_RAM_23 => X"4D308D468A15721026228A905488C2A6015A02518012B2090E14840AD5404814",
            INIT_RAM_24 => X"0410A915696A20E42A5540A8040881482450018F3131DEB900033D0159AA2320",
            INIT_RAM_25 => X"A1C8214034767F874341470000802AA8E00605C202202584A5510546A10A1081",
            INIT_RAM_26 => X"030500408E08900A0B402256C44010850412900A013328BFD8B15454048D2852",
            INIT_RAM_27 => X"39404252913E04F912022186442C329BA60040808780218F25508858D6252A21",
            INIT_RAM_28 => X"889600C6A1841A186810100200654322086184860108104D8690C961B0466A04",
            INIT_RAM_29 => X"4822A14C480150956066244102589401687CC000D8393021CC511010968121C2",
            INIT_RAM_2A => X"607BC80528850F46D5A2AD51210AD120E228180210881250A428020583440409",
            INIT_RAM_2B => X"223234E4C202D88184190342A4F33503F19CAC07706ABDA0886A51034BA9585B",
            INIT_RAM_2C => X"54841441E128521CA548043516962512A264350A92505254A22200B490128140",
            INIT_RAM_2D => X"010020520811010052C2100BB1041B12AA1111091420822A0096310444814095",
            INIT_RAM_2E => X"2B805165409A8B6C13844A0050181830810088D8180002204448A048101AA990",
            INIT_RAM_2F => X"3C0D49C0500057A5125410D80612402209140209268D625C024940504C20101A",
            INIT_RAM_30 => X"18355488B545AA262E902913494A4A654A0410B5D5824A98F6A501CC7B50B6EB",
            INIT_RAM_31 => X"06DEC10D5604A5CF0175A0090B10D0FED8727046004100C611A41184AC671A01",
            INIT_RAM_32 => X"0AD00EF7ACBA80D8823AC92053549975B128031684920F2B124B42A2B0AD30A0",
            INIT_RAM_33 => X"10015541228208465B12840540340202202025807949221429A8753F1A279501",
            INIT_RAM_34 => X"8285440264881B06B60C92FB00200026A2005A00200AA00E2884341049001B90",
            INIT_RAM_35 => X"9A880004155482AA010841041000011100900008042210022A8BC80000800304",
            INIT_RAM_36 => X"640023D83046C1502A896A1AA44102D149C038D1130A24084012993890A89000",
            INIT_RAM_37 => X"84A34C500979389A580C440E00B828F1A0B735AA1205177553D2085702421505",
            INIT_RAM_38 => X"802505C54D1C8110010489912348802004091092AA12502A33A10AC0AAB04A9B",
            INIT_RAM_39 => X"E2603881E04000EE922AA412602C1F515464ADEFACAF4A045F556F4BDBEB014A",
            INIT_RAM_3A => X"54934E7821AB444056A2AA8C8247F22624305F6B8B21FE538D9416480C46F525",
            INIT_RAM_3B => X"C8650001931B649316A0FEA1CAD50264C8593CE68428A77669A762B664C94234",
            INIT_RAM_3C => X"2C9A84641FDA6A351D2866762840321EA8E90A5943147A97F202262369618156",
            INIT_RAM_3D => X"C9226341547AA0AA600C60ADFABF9652C36935B101BA224470C319009F93FEC0",
            INIT_RAM_3E => X"0525844B436227A448A7646AA448DA495E3B34ED21A3AAE319134C95042632DC",
            INIT_RAM_3F => X"4B5082A64A595C54221E2C4B5A41441075369B692DFE943114B58099FE8B73D4"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"D31B696680BF2C34F4F4C1D11E8C6D0CEEB6A0D04AB292125A57A21825D11A09",
            INIT_RAM_01 => X"3D862BA7973B6B976ADFEAE9A5B7F850105454545400E770100E1D8A1641AB65",
            INIT_RAM_02 => X"9821C10600FBBFBBA3D5AA69F2E45EE9F816BB6B11F82A46DDDA6FA1E3FDB465",
            INIT_RAM_03 => X"057FDD6815A75C23EB7CFD5D54732E5337CB74BDFA1B15E20D5F26997DB0A3B3",
            INIT_RAM_04 => X"AB5D3AF6B5875BBEB4FD1D3FDDBAEDD6B4AFF7F3A1B7DDF77534093E9234C802",
            INIT_RAM_05 => X"25A7AEFFDCE3673B56FBB2294D2BD418A0768127E9FCF6FEEB4BCADD6EAB8C6E",
            INIT_RAM_06 => X"092C20480934440E3DBBF0A030809E0906A753353B00A2005BBD4EEA7FB9FA70",
            INIT_RAM_07 => X"C83EACD0058FAA789DA401440AFAC0034508B0F1EFF5A35D80918C049A18A434",
            INIT_RAM_08 => X"A000915229829D281679013412A24204AE38780941E054A1010888A05DFBD3C4",
            INIT_RAM_09 => X"041350C020008B32392281000022400A08A88191C65D0D60290C031ABAB3FEE0",
            INIT_RAM_0A => X"3B65C5800C93B15FFE35FDB49806784804108A76213B0239A5008A20010C22C2",
            INIT_RAM_0B => X"189A63A4CD0B9A0324214444191522668AB29930CEE049B465E1011DC20A5142",
            INIT_RAM_0C => X"A23A09592058414428353F17C8C7B151E14A150200544045050090C677D8A38E",
            INIT_RAM_0D => X"2C499444006CFA9918A66D19C94A6032714E1B2D0DD4D29294ACABA45274D187",
            INIT_RAM_0E => X"334BBA145106519D2B12631880009B82EF33FFF7D2E1F9BD0AD3AE8537E42595",
            INIT_RAM_0F => X"80B2959E02285191AE5930810430010CAA210D15423C755848E271FEF8F9C0CB",
            INIT_RAM_10 => X"566582020665A1900A52D04A208032953012811845042048848920B5A8A101C2",
            INIT_RAM_11 => X"D0C3449A33006AB23B109CD004911C0C08922A8BB5229026E18D51A439086026",
            INIT_RAM_12 => X"28018C04108E10C729045D2A4283B85E19147482459E59467091546B2C9AEEA4",
            INIT_RAM_13 => X"922884492D81082F5E198258E2609222098995666780213300471A68182319C6",
            INIT_RAM_14 => X"C5AC8232E5C2C38A4BFFC4A9472522D499116B411D036002894457232613FB64",
            INIT_RAM_15 => X"26ADAF788DC186D01168008004FCF76D451EC3CD60914710137CC4020CBA6317",
            INIT_RAM_16 => X"41703F048EAA104A79493E0A443080A4A2970B9813E7ABBCA00B60AEE57417DD",
            INIT_RAM_17 => X"995161102C2C210506555CA14455772A02FB501510042084225631D81D973BE8",
            INIT_RAM_18 => X"0D09977EDA5311CE22360D837B60286D28F4028789C23285AC914001012150D0",
            INIT_RAM_19 => X"64154CB00E661462E4C6994128A208CCAAA200184142C2E4008AC8596930D03B",
            INIT_RAM_1A => X"0306CB361FE49385B284593201729A690C1CA58C61105000C618B2B40431C8BA",
            INIT_RAM_1B => X"B8B385866D8F3E2AAD23CE885C806EC95DC2208AA5F4444432A4D933820B0803",
            INIT_RAM_1C => X"84508A802243100830CCE45421031C506C50A804B117C26792805318C311E458",
            INIT_RAM_1D => X"6DFE81B53CCAB560A4431BA55DB5CD28CA16321C0348312CE11001B489DE4431",
            INIT_RAM_1E => X"28D1E9E005E5424617A4826915BBFDA5430831B502A0A28082F84B5CF210EC46",
            INIT_RAM_1F => X"81C0235546440AABAF588D9CB3DF6CB3D9F519290BE95557FFDDA40EFBA88414",
            INIT_RAM_20 => X"27F84632542BFBEEEBA038D2118C2BE2226BAEA0A084529402408960100B5812",
            INIT_RAM_21 => X"32AAFFF8A5F8420FBC514A528126300582998002D2B7F12A949613FE18E39294",
            INIT_RAM_22 => X"0484E88F7F5F12220131E491216042DE4436118E50B16282608618955DD77204",
            INIT_RAM_23 => X"19B8CC4603D9EF13468028A15122EA181EBFD07A8139531D0230C0D071DCC383",
            INIT_RAM_24 => X"30508920F028062162C40A211CA8038875181882A930F7E787218B307DFC01C0",
            INIT_RAM_25 => X"C171040874303F0F034544000084000082130582026A84D4AD43845028C58F3E",
            INIT_RAM_26 => X"CB24A22A541C4A4B09283256CF156006102B00A8003E175CFA81DC8404818042",
            INIT_RAM_27 => X"D424421E1DED37B5D2832180042CA0960CF1FEFF31117375DD42A117ADEB6820",
            INIT_RAM_28 => X"2CEB128A25008A500E18B4809D544A224940C704210C0C0E06F1B562F0C6A606",
            INIT_RAM_29 => X"02498D87842078112403C249204190483DFDD288483B3236F811F348514610C6",
            INIT_RAM_2A => X"B84842641C058922A1822CC989A2D802C02233C5AD1C3A78F4DF2A4483408480",
            INIT_RAM_2B => X"57EABA5FD08C5FE3A137C7517F437E00372C4771BC9E49C2284011070C8F684A",
            INIT_RAM_2C => X"B1AD3D13CE729019CE5110CA76A1CA440030141836D4D4C211E167A9B4B613D2",
            INIT_RAM_2D => X"18C390D22009904B8F98838516DBF10675CCB492EAD3FDD433BA0EE3C2375BB0",
            INIT_RAM_2E => X"4357D26814582B8C6145FA287BC8EDBCA4425EF29AA119068005220809A5B4A5",
            INIT_RAM_2F => X"890AE4C911401B5CFD61205AA40210100B404304007191340D3E164007A4C361",
            INIT_RAM_30 => X"9836D3CAB4C0F91B1CCC004D813091B32212088A5C5A088E631C644530C49A44",
            INIT_RAM_31 => X"033C6826D20393ED10301910E1D86834821E1173804884210C40134002110440",
            INIT_RAM_32 => X"0A152226C20C520E488860C8458426B4F00929DB63641200D04088881DA6DD89",
            INIT_RAM_33 => X"4A086C3392C20103A267204CFFC2FDC0A2A2812A1262C9808C29145B0E9B6028",
            INIT_RAM_34 => X"1D0C4C12128A0A51AD57DBE0F69772CC51C71CC32C60282A5B651127B3F15919",
            INIT_RAM_35 => X"B1471CB121453E802A5A642AAAAA943AC9D45410402694402098176DEC566D00",
            INIT_RAM_36 => X"32FB47A07FBECFC4B86D3353F458600A11B2340BB099CEDA3398D4968049D555",
            INIT_RAM_37 => X"CF81B40D5DED368E924D83443210A0E508322102111934263DE704231EE3163D",
            INIT_RAM_38 => X"540172182024A950C065A5BD47FC9C217F081003BCB30C780C101EE1BCB0F86C",
            INIT_RAM_39 => X"10190B08420004447458500013238A32CA1008DB1A963194B630470191A89A25",
            INIT_RAM_3A => X"8225014804CDD7141AEF06218DFE630030094518C6D87C73DC12DE0D02412291",
            INIT_RAM_3B => X"1A98F104CD0D936405880C64A983003340064C7383001C0836D81831BA231105",
            INIT_RAM_3C => X"21761033842C201400C0330188E5B5E3009918380014318D9DA4C1CDC31E4AF1",
            INIT_RAM_3D => X"3259109209318C1298221A0B19624184B0B2C18E04C2C90BDCC0410004889226",
            INIT_RAM_3E => X"309B391380F8131B04D0C2205D242CB35F09122494303204866CED68C10B188C",
            INIT_RAM_3F => X"D45420AA42DB4B0CCA012F31CBC55C4403DB6D9648D98B4E715AD40C6E62399B"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"00995682102F2D2A6036164840850A0201B73A425C4490961364CAD020E8DA1B",
            INIT_RAM_01 => X"6CC31850069A48044194430C30548E63362776633621E7B3637F1F10927E5C1D",
            INIT_RAM_02 => X"01044B131802328980810C1427A4119412102C49926820039D5F07515041A524",
            INIT_RAM_03 => X"5A002BCD40F82F9E577DA9F77DFA8E79DA62FA28210A50E8009814267950A383",
            INIT_RAM_04 => X"4514423A98CD809B06680C428CD2669319AC0909977A7D5D7D57D421C2B3FDFD",
            INIT_RAM_05 => X"81D1C8046C25662A033B188B1048F29D50182002800AD22C3508E04443482643",
            INIT_RAM_06 => X"310D8C700870A1FF49824D204B2C07490F0F4409444D000C1F8C14347519D010",
            INIT_RAM_07 => X"4A001209AC350057A46C92A3955606C4282049ACB8AF440805A9BA9515A88C50",
            INIT_RAM_08 => X"52B22A2C46394A8405560814152B82909860794D8151080484E121010A74E484",
            INIT_RAM_09 => X"70062E8BB37776D87826E2C04264498B9B3B19C2AD89001E9253A042E0668D23",
            INIT_RAM_0A => X"2EBAC1BF7284F00AA84219271064D39DACC31A88694438114A8201DA1211C048",
            INIT_RAM_0B => X"C08A00F0481F996B00031025082DC07A132B88105B8472A8748608000C0A4203",
            INIT_RAM_0C => X"687ADBAD049B4A74046A1730429F2181C083E999C688D9DDC68781C6E9D15C30",
            INIT_RAM_0D => X"204809A50C810501915EAD6B50226A1A249A944AE22CCAF5AD6B0A11A6E991D3",
            INIT_RAM_0E => X"F00E001116440100270528C10196B60D0A000000092C0E021BC3C099E5E22512",
            INIT_RAM_0F => X"48C1191C680702282004431A018219EC44522D8007162088952C91C282885A37",
            INIT_RAM_10 => X"0007009280070307246BF40A3816748162E527298F7CB180C08B05112B3A894E",
            INIT_RAM_11 => X"041072D27268D5CC486C10A0009114556408C51400787402E08D43203E21A906",
            INIT_RAM_12 => X"2B09797EF782949C8C40A02D0082342E001C01C54230C31E6046885368188E30",
            INIT_RAM_13 => X"69C04C64920C63C84C26689545C52A88E4F94D4C453446A4578A234814A56B5A",
            INIT_RAM_14 => X"CAD280A88309042012000F0C4847FA4C78B99C847646A4CEDC41DB1304B116DB",
            INIT_RAM_15 => X"4624808770FF39334122A81A72C0BA4D401B1EBB8C500644000C48A81243AD15",
            INIT_RAM_16 => X"CC82C2404B114320504489012838708B282078C18EA501A93075C2311A882822",
            INIT_RAM_17 => X"22001834D0D0C600802A8B52A3A0221111024104011106F3C68DF22122141141",
            INIT_RAM_18 => X"2200022BB55CA90933C9D266D1E0B920200805427220E8AC60802CACA246A300",
            INIT_RAM_19 => X"9D4279431181C186A24460AA0212971501AEBBD35E3232009A9503106903A344",
            INIT_RAM_1A => X"2C45A06D8D210F9B4D0A0054C020D00B2F02198846EE03F098600D4B9B080101",
            INIT_RAM_1B => X"39540350907280000180C5240A4482180A03C0004005DDDD2D22B44D2CB6558D",
            INIT_RAM_1C => X"900F81BE0D865C39E0122908C604000E23081E6735801200641D0C630190A40D",
            INIT_RAM_1D => X"900004002883A80291A090180A230301EC0463589C27CEA03AE13920347FB865",
            INIT_RAM_1E => X"8102043C4140980039006D0105B9460A458453D0A84FD99B1801800020329344",
            INIT_RAM_1F => X"66C06C00003964000018004418618618600008708003C820820008E000046600",
            INIT_RAM_20 => X"CD118C6001940411555AE8D084211408602AAE85A350225483063CE0200001C4",
            INIT_RAM_21 => X"9C5145148AAA85B20A209800500220C1000D0322FCC1704E0D08668861860008",
            INIT_RAM_22 => X"610003001400790809C8E40816002904021908400140600882082002F22009FC",
            INIT_RAM_23 => X"1148281422B146B1003BBB00DC0C0EB420140680045004AC665E1C1038407820",
            INIT_RAM_24 => X"C01D2F81A6F3BC0142840120728E0483078230A051B3EFF738477A0DDC8844A7",
            INIT_RAM_25 => X"91720088F4347F8F870527004AE299EFA53EB5739B082F07C9F87FE6223060C1",
            INIT_RAM_26 => X"2030118200C040C52501650880608B1881804221020BDD9A8C78605846B0406A",
            INIT_RAM_27 => X"AB4D5B75864999267D8A2D14F68CA08628AD54AA61840400000A302CA529480D",
            INIT_RAM_28 => X"1BE1A6D5CDA114D834D9220C567B9B44DB60CBB4D161974732A031C3F40C8AEC",
            INIT_RAM_29 => X"E48023E86803551861F434430182AE1B482A22B890826CA0019800443C20CD9C",
            INIT_RAM_2A => X"C05CEF2781028A0A360890640A299282A40B62B3188A1754AE00EBC10812060C",
            INIT_RAM_2B => X"300516A0C05C800580802B0A80250B81E7CE6B15DCA3444AB18B123011D443B5",
            INIT_RAM_2C => X"1D29BDCA8A5016316A43109CF6039C30BA5A30D264849491820A892926A48515",
            INIT_RAM_2D => X"6B56A9C84283854250028618000062140025416A00A0888B251A8014550A0524",
            INIT_RAM_2E => X"0310656072D8C1CA4C34414056BA1A100180C05848AB6AB228800D09B880C003",
            INIT_RAM_2F => X"C99E62C8DD8C81DEC966A706D6108136391088992C34381029306488D6874489",
            INIT_RAM_30 => X"4042631E8460C08990C4A1C49A39989928009A08E05A48843118C46430CEC800",
            INIT_RAM_31 => X"C3B06846D04B01009431989CE18625B0D2C630033648A52960C0936022394678",
            INIT_RAM_32 => X"6E062770E62E02CC489870CC0D8425BCC00B318163641230E08084CECB32CB09",
            INIT_RAM_33 => X"44A74051448B4C1461E0B1A0631263113BB3313B32E6F1D899B9064B8E59248C",
            INIT_RAM_34 => X"FFB475263410C80F0C4492E3189C1288AE180C184001844C1E60A5E371BB0802",
            INIT_RAM_35 => X"2AB86180170818B9381105E79E79E009A856722DB60911E453E3FC9420CC903F",
            INIT_RAM_36 => X"16026B2018065F9C888262822D698C482AB8CE5411BD835AD6A0448454384675",
            INIT_RAM_37 => X"C271B8CF0E0F47A083039654E4328227120A63388A70C860780384284632C701",
            INIT_RAM_38 => X"080005F80480A34280EDBCB77FCDEEFE373A2181AA70193B6D4A6400C383266E",
            INIT_RAM_39 => X"C7BC1F2CEB23210064828ED0BB2B0000001008DB1DA635ED3630470191D12490",
            INIT_RAM_3A => X"80252841CD8B142374A2E30B30C5DE428D580F3186D8C0DAC531221C264B704B",
            INIT_RAM_3B => X"53CA621CEC6C9B247500EC7520C1B4BB1B1304212B8AD94896584865906A166F",
            INIT_RAM_3C => X"496495BB8C668164BA6219849B3BA93EEF8BF3937881B1CDD933C840693EDE63",
            INIT_RAM_3D => X"B2C935B683B1810792221209903241449D96512540C3C0201E4A60670DE1B26C",
            INIT_RAM_3E => X"E84B391356E8431BC3B6E0DC1D0D6DB3544CD9B2CC2E2490224D85F853594C8C",
            INIT_RAM_3F => X"9820B4AFF3FFFE19EF7E7A4A5E91F9B6F94B2DB6C8CB93989918E12C6C2610D1"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"259110C58840180222366049BD82008A21240C7105199B3201423DD804A25002",
            INIT_RAM_01 => X"9134C44AA1259758B4690471C4C8148C8DDDDC88C981CEA5A8DD9B331301A288",
            INIT_RAM_02 => X"A4D21244450D8946766A71904C59A0228445C0A26607D5E43E10B82623220B89",
            INIT_RAM_03 => X"8D72236DE577D8E88A2F8B28088DD188251D09128600E402B0015A4A82030C10",
            INIT_RAM_04 => X"AC88200000301F203892D02110048020410329DCB77F7D5F5FD68A21C2BC2A88",
            INIT_RAM_05 => X"104A240290848114400087243C800A829601D5842C0700D15A6008198CA76B8C",
            INIT_RAM_06 => X"52C8B344DA22000852A4A64D9B6CC1840112384380820122840120CA82220D40",
            INIT_RAM_07 => X"031459A4B60050D6D73602892505025832A24228200D50004284924A54A80602",
            INIT_RAM_08 => X"58D8662CC6610AD01DD4259B38760FC0C9A1870A20040E08A0B414510000D8A4",
            INIT_RAM_09 => X"1A022C2CE0013241249130088D11260E4666C468248032C3296D0CB12722954D",
            INIT_RAM_0A => X"28A2090B0A5892A028AA82491310010246A845A913D4851000D2218CB9B00003",
            INIT_RAM_0B => X"60C481520082012417B4E10A000711114ECEC6A362134080C09081B3211828A0",
            INIT_RAM_0C => X"411112A48D09C49C010290554D728AA8162492113372722734B44C64A9735C10",
            INIT_RAM_0D => X"902CC228E1100000935AB5AD64010503208B009ADAA84B1CE7380D40A4A9055A",
            INIT_RAM_0E => X"642C00188092A0A03260442106F100D040A62AA2809880E804491222200A424C",
            INIT_RAM_0F => X"5214C33048840E6E7932C84C865423140084150282468AC83323908305064780",
            INIT_RAM_10 => X"B0B11D8000B1165C844241B4C65826648908590D659EAC363888C9864EC6629B",
            INIT_RAM_11 => X"332D9A428A625109042362A99A2900E0C76B6B810210299926C2C99A224D4444",
            INIT_RAM_12 => X"BE03190618C3118C00A008912BB040ECED09826120102062DB5B5C5246C41C13",
            INIT_RAM_13 => X"0419140000040099310CF5E54C0EC46580B2669108033A83240A612CA5C5AD6B",
            INIT_RAM_14 => X"1B566CC8896430C68400908098400499B20D088D931293131085347250000000",
            INIT_RAM_15 => X"029329CCA9A1000CDA4446409C800C923600500028DC8333000C8E4EC30C2108",
            INIT_RAM_16 => X"9288003B324F68E5011C810D4613019920F8888448300100C0011EC000080002",
            INIT_RAM_17 => X"E604008B52521080D9AAA14289AA28C46E098CB2DDE6010191654624E248D011",
            INIT_RAM_18 => X"90866282022081082300C02000C886134408151200086CC630C426060212A928",
            INIT_RAM_19 => X"08E83348F090281131656EBCD143313615330120608707081A3123640488A9C4",
            INIT_RAM_1A => X"A0401A013048C64900D4D22488004931A3A95510D885A480A104014980421241",
            INIT_RAM_1B => X"8354083601084022209291B1A2531108200211800A022222248A030124924600",
            INIT_RAM_1C => X"D108D5841C82611820899802108269ABB802188CD700344D5F42000004DA36AD",
            INIT_RAM_1D => X"494038CDA69A2A9093203018AAE23365A10C02480A90213126A00726445AA826",
            INIT_RAM_1E => X"891226A886463424101A70504730043041941B6A75000CC6640C2CA0231A4844",
            INIT_RAM_1F => X"35C05155578288AAB20022235441041042004424E01100000028021100026644",
            INIT_RAM_20 => X"0002108406C00000001C320000004002484A2C8122004A85200008CABC0D695E",
            INIT_RAM_21 => X"2800000150047A40410C0B1040840090804819CB418044374E01000104104001",
            INIT_RAM_22 => X"B05114401080100083049CEC5940B280909042100009240000000002C0000402",
            INIT_RAM_23 => X"1301383C1EB34A89A14444D6269111D80010000410100008C2110A2552234458",
            INIT_RAM_24 => X"C09A4C5AA2244C01C18280F01481412486204430502063F558454D825800110A",
            INIT_RAM_25 => X"1044C02878703F0F0F07650008D211B104228B04E399042619C4004B74102040",
            INIT_RAM_26 => X"642144D2A9A3148828510010959541C8920A0D22078ED587FF28422040905009",
            INIT_RAM_27 => X"00002B0008922248808615191418738249AD54AA410200000002200084213511",
            INIT_RAM_28 => X"40C102C02588025804189AC150604B024160C2D488A14920900C13602276B326",
            INIT_RAM_29 => X"01965925021C0659B012816180866A04208AA1DC6BA18A4552315CF1300C6602",
            INIT_RAM_2A => X"40508040200481404410215204028090090026A5290896010CAA1E66BA620C04",
            INIT_RAM_2B => X"150512AA5B592158B682912A8003700229DD76B397B7D81004205480210460B1",
            INIT_RAM_2C => X"1210962810035B02202990948252958ACD914E2100080A18CE9E841202C04D2D",
            INIT_RAM_2D => X"AD62ED400940A0A4402148404020261800234F6400000089C400C44D2D683402",
            INIT_RAM_2E => X"214548A58A49152084120194042C0A12522340435A318CC7002C910ACD008DB1",
            INIT_RAM_2F => X"1210B00E2260F01482CCB0D512DB2937282E2E42015329ADB20B53A224B6401A",
            INIT_RAM_30 => X"362C888B688A2CD2E9693C2965AD2D2A91C9B650B6A699294AD698860D699611",
            INIT_RAM_31 => X"120907102088C298198C431214774401661425CA5448C64202B913B995A2084C",
            INIT_RAM_32 => X"1199E45C9D89CE6B9816CCB16A2B580A239424765A8315850E3961B3304CB056",
            INIT_RAM_33 => X"0407C2C943B34D1B20C9322000340014664CC0142094856396671D90E1234BA2",
            INIT_RAM_34 => X"344CCD8A33C509610509242DBD825129AE0809041064D59428A2A43018000CC6",
            INIT_RAM_35 => X"EEB820C09DE2B6444D456634D34D0193249DDACDB63148418418124948C44B02",
            INIT_RAM_36 => X"4AA4B0011552DA6625BBA686AA69A0D3529926C1200A2D6B5AD980080A0C8CCA",
            INIT_RAM_37 => X"32440223EF432188726B2226131B84B184E331850DF009B4895B06C4A946CC2B",
            INIT_RAM_38 => X"245488320484C58C84CEDCF5DECC8E69B6148821AB3089B520238590E9AC2500",
            INIT_RAM_39 => X"0089966C932018112185812A2C11409C301A92004180804C008090A824011452",
            INIT_RAM_3A => X"2048214812992C9D919212521044421207108B2C2490816722C80268906A5802",
            INIT_RAM_3B => X"5B803580650DBB6C258F052E3048811941210B4AC10B099826988018B30B3B03",
            INIT_RAM_3C => X"B3660819C003250C8026190804314B6032815A0DD08814A489002E82690E2E30",
            INIT_RAM_3D => X"16D8A120228400422515A51024049249012492CD08059020044CC20240080216",
            INIT_RAM_3E => X"025243246085004090188805028D4105200D9B165A040010888945A20A121523",
            INIT_RAM_3F => X"980081385E492F89A020AC842B3968B009924820921202101010984C4934A522"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0836FFEF41004AFFDD07C28B29A99A5131A518A410513E2680A0567CB2843400",
            INIT_RAM_01 => X"00080000000000000000000200000262622623333322CE8BFCCDBB9E02820808",
            INIT_RAM_02 => X"0000000000000000000002200000044108020000000000001C0F001010000000",
            INIT_RAM_03 => X"0F5A81E7457578B5A220768022880A4000000000000000000000000000000000",
            INIT_RAM_04 => X"100204004200204041002200220110080210D74BDE4F1D580A2B5FD6A5774A02",
            INIT_RAM_05 => X"0000014001400880080440008010012000A00040028009000010012010100010",
            INIT_RAM_06 => X"581A69ED6C6991019AC6827B114D958B6202F736A6D8404020420101004400A2",
            INIT_RAM_07 => X"F6DB67B260CD7E080880A40208796933E4D1ABDFBEB48AEE28C2C327746C8D5D",
            INIT_RAM_08 => X"018104D89DDEE5D3B758A298F22E5A05CCBE84C25741F1534F26761AAF153525",
            INIT_RAM_09 => X"1367B13AB58BB6E586E1256819B192D6092E48CD36C8B05FDEC45456B2279F58",
            INIT_RAM_0A => X"EFBDF021F17136ABE9EBD2493C5CF2D4AD252498824C4CC3F0359628E9F60D2E",
            INIT_RAM_0B => X"2D10B54896C86590CCDDDCD8664DB53122560A68A249EF41420A52A814ACE416",
            INIT_RAM_0C => X"4014C0F23187F4D7817EE858345251AC19345A11A7C176675B5A11F03D5964D3",
            INIT_RAM_0D => X"D6B33A37D3360A23F963B7AD6EF0D58C67943ECF97796E56B5AC5941A26880B2",
            INIT_RAM_0E => X"80B9FFE0FAEBFEEA60C3931A790EC93830D0541C76524DC07E6D49220A0BC870",
            INIT_RAM_0F => X"64683A53BE5BA72309FC4D6CDC0AC583332942E81DF9A525B9108A3DB8B22099",
            INIT_RAM_10 => X"4F0E6250AF0E5864C1F7BD41837ACB9A0C62244F0DB7E68B45C232FAB6E5338B",
            INIT_RAM_11 => X"88ABDB2F4CB0F8CD8468CBA2C4038E7E48CE49A0C06A86C5390A6BD4AC93928D",
            INIT_RAM_12 => X"5EF1AEF95ADB68D7C2B106E9F4C8020D14A8550DB0D36C9307724DD120210D0A",
            INIT_RAM_13 => X"6885BEDB6DF2734E9244440347131B1C7AC0CF2190110EC4DC5A30DEAC3DAD6B",
            INIT_RAM_14 => X"0D7B015F1838EB89955A634289CFFB2081437B224187C9B9A0BB921E589F56DB",
            INIT_RAM_15 => X"8F501086F20646F92599D572093E34D820C538409D713380E6AB3381AE3494A2",
            INIT_RAM_16 => X"0C8E0044832DCE318296C1B9B99AD5FB310E1EF17E8FD4415EF769427133430C",
            INIT_RAM_17 => X"C1F2D2C88B0B1ADAC8D428A4020F8F4CC45408C308C65E9F408A0262263C65E2",
            INIT_RAM_18 => X"405728F324B2C0C623C964890E0770DCB7F2080D4C06980885B2C8909458CD6D",
            INIT_RAM_19 => X"E6AC01C4158DA90A4D8BDA20FB4D0A6874C03A8A81804059645314CA1A6544CC",
            INIT_RAM_1A => X"9429249240303A6D92392C4936843753F27FFA570F70EF4518A35884D810B05E",
            INIT_RAM_1B => X"418C5B496E705499984D7E54ED1A112EA837FA7550F888896D4B2493145BAC30",
            INIT_RAM_1C => X"6CB72A424588AE650D1003AB58DF3CBAEBA3F9168CEBCBE5B263ACA42867D952",
            INIT_RAM_1D => X"261FD37241656BE7DC36976BAFDAED9605ABC4872127CE5EAF6242496762D88A",
            INIT_RAM_1E => X"C993266EF9B3B498B5C7DF9C2C4755F42856842F6790D402ADFE3EA99C44132B",
            INIT_RAM_1F => X"8440A55541EFA62233879999D75D75D75FFF7267DFF2AFBEFBE74D35DDD98B64",
            INIT_RAM_20 => X"4756B5ADA87FF7DF7DE2113FFFFFF54F8594517F5DBFBDFBFDFB2F03EC0D6BC6",
            INIT_RAM_21 => X"C5F7DF7E7FE6DD2B2CB2DFFDDFD9E7E845F73A752DBDA24933F9A3A9A69A6D7B",
            INIT_RAM_22 => X"88EDB6DAC2AA76CDEBF753AFD2DFA5B7AD76B5ADAEAADD745D75D76B0BBBBC00",
            INIT_RAM_23 => X"E8B5E3B34468B1A63C66661C70C98882F540EE5DFBCEA7E258DCFBAFD1FF62C5",
            INIT_RAM_24 => X"B59349E206F452FE3638FD1FA775561EA59E8F6D7A6BBD6C7DC884F823AEEA5F",
            INIT_RAM_25 => X"EAA3FFD8F0F01F078B870105429080F7C11DA6E6E3E9AC64C17606C1477EFDFB",
            INIT_RAM_26 => X"5A5F417DEC3BB596F6D7E6FF332BD3D36874E3DF019E38BDAB7B5B8FEB4A8EB4",
            INIT_RAM_27 => X"F78DBEFFEA921B6CCB77DF68FD7BEFA13CB377BB8A66E6BEBFEDFEB2B5AD4F9D",
            INIT_RAM_28 => X"0CDE7DEB5BC2A5BD41FD533C63E6B78DBEF5EEBD3EFAE0B04BA50BF82A8F55F5",
            INIT_RAM_29 => X"D56E2B755B4FAC8B06BAAD8C35119F63A283C60175515D5D7D5B4411F28EF739",
            INIT_RAM_2A => X"A0610C8BD9EB578DDFCFFE4BF1FF336DFEFFD0442160EE815DAFE30F55C4E4DE",
            INIT_RAM_2B => X"D8286B05676080AACAC155EC00168401E18DEED0A5BD5B8FF0FDEE0F8E1AB134",
            INIT_RAM_2C => X"594B634E8FD56679FE8C958C7B58C64B08C6FD74ADADAFB6B141B1716DAD6283",
            INIT_RAM_2D => X"39C7B27F9562C75B6D1EB3673D96B3759E58A0D53386EEEEF975B32A8382C16F",
            INIT_RAM_2E => X"B5A862364B6E851A4BCF7F22DAC7F7C1491475B77563198E5F72C9F78B5BB24F",
            INIT_RAM_2F => X"091846027770F1061A4CCFFD9FEE494A2FF73E3268399A9FE588EA3330642B65",
            INIT_RAM_30 => X"557C0899AA4A21C9CC07EFC08690809895AB770A7277BCE419487A2290E78F04",
            INIT_RAM_31 => X"191D3EB06B8959C88F8A4D1C345F2B8040B196604C4C6301E07B02BB5099640A",
            INIT_RAM_32 => X"CABDD0167CC5ED80F5C38E69E621399E69C7349E39CF93F4ED14F63BB32C7349",
            INIT_RAM_33 => X"7CF89C1EA76061B06C064B395ACB5AE266666A5E946230974C06A10144B101D4",
            INIT_RAM_34 => X"00BF6F5B4BA75CF042A9A4B939AB8D3CB269A861A6D897D9AE9AC8CB65B3F336",
            INIT_RAM_35 => X"BAC9A6DA2CD2F7A665A5DDA69A698B7733B4CB89A6E2789AD07C009EF52B24FC",
            INIT_RAM_36 => X"A306DB1D54CBA040F01CD0E4DC04152CE6E5A120CD3D396F5AD7A3F9E337B5DA",
            INIT_RAM_37 => X"74CC1A2467E3F1D85498088DDF57B9EB7126EF7059E41B2C1B49AD4888713455",
            INIT_RAM_38 => X"BB16A100B657874D28149D977E69AAA72640000A6909A31C531D299A3FFA4D06",
            INIT_RAM_39 => X"982240121CBBB3CE60303EFB2862746D96B2D8D21956258AA432C72D218238FB",
            INIT_RAM_3A => X"0B009DAFC0C98E0051C6E63349F6664948C34795324245D68A624BCAD4F1236B",
            INIT_RAM_3B => X"7EC26AFE89E922499B760C665CA078A26282E3019AA61B02820A0B511627A788",
            INIT_RAM_3C => X"602DF7A2E309B4C4425180A8AB21437077C33D09BA7BB18D9B481010C38A3A79",
            INIT_RAM_3D => X"260B848689B191568452844A81501864A4105881A85005968178AFF8646C8D0D",
            INIT_RAM_3E => X"68C981124C455B13053002DC58B20C31A0E040228852C5CAF4A037A2E8484D8E",
            INIT_RAM_3F => X"3800103DCA4B3FA20540FA94AEEBD262F301051458C2210CCAC6138520601868"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"F7D92100BEFF8C007C804E11C00A000000251EA0105D02A00002975900F85B89",
            INIT_RAM_01 => X"FFF7FFFFFFFFFFFFFFFFFFFDFFFFCCCCCCC8CCCC8CC3848E5A3812AE80022A0C",
            INIT_RAM_02 => X"FFFFFFFFFFFFFFFFFFFFFDDFFFFFFBBEF7FDFFFFFFFFFFFFE3F0FFEFEFFFFFFF",
            INIT_RAM_03 => X"F02DD612BA8A808A22282A88022A082BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
            INIT_RAM_04 => X"EFFDFBFFBDFFDFBFBEFFDDFFDDFEEFF7FDEE596D96480A08222A2A82A2983FF7",
            INIT_RAM_05 => X"FFFFFEBFFEBFF77FF7FBBFFF7FEFFEDFFF5FFFBFFD7FF6FFFFEFFEDFEFEFFFEF",
            INIT_RAM_06 => X"63ECAC500032E0AD1284834B1240050821F355584087BFBFDFBDFEFEFFBBFF5C",
            INIT_RAM_07 => X"485961A024000659A46C0AA28D01001D780898633017908044041A4640888412",
            INIT_RAM_08 => X"F0D032664A570E008A0828A22C57855051447DC2821104050171114000341C20",
            INIT_RAM_09 => X"600411A3211C84813095404B0F552E8F145DD8C9A9098A36D95A228CE4669C5F",
            INIT_RAM_0A => X"4C30111550152000280012491B108211074844C91264B55010C0823E0BA10007",
            INIT_RAM_0B => X"A0028100208B09021E03556100231229578F8E81731450882694842AA90128A1",
            INIT_RAM_0C => X"6F98D2001811E69ED040510025EB3128D2A7A38804989BBBC485017481AC2020",
            INIT_RAM_0D => X"900602A1EF70000028200C00042205040618404104420A1084200B400481150B",
            INIT_RAM_0E => X"900F505B9282B4AA156D7AD00142240506904010402405803D08DCAAC162515E",
            INIT_RAM_0F => X"4080021AB2090771440A22160C840100445200028850AA48F7A7D0E864614472",
            INIT_RAM_10 => X"000028A00000134EA0C0010AD80E12C129C20A0C2F267000108180940D5CEEDD",
            INIT_RAM_11 => X"2208AA0261288001440A0204118900E0E22A9414280530108C41491120002586",
            INIT_RAM_12 => X"142821282508041088A0A0B52199FDF6450428E90A20E2286154A08247DEF622",
            INIT_RAM_13 => X"69C1DC76DB0863144CAAA9F0A83E2889C8DACCCD57A444A04A85420A00080000",
            INIT_RAM_14 => X"F9D2FF68890DB6F78CAA0708DC4000045AB1CE18AD44177754C03903101D76DB",
            INIT_RAM_15 => X"0224A84050D22D8F0003374A7669A693BBB41440084EEE7BE2ACC0F7DB662901",
            INIT_RAM_16 => X"54482831525848010040A11D007210BF2804FAA0729554B064554068C4600618",
            INIT_RAM_17 => X"7710503258D88400D56A834AA2A0A0FFFFA2EEBAEEBFC17ACFCC37A57A4AB400",
            INIT_RAM_18 => X"9E8D5A0224688885106D5B44812A218805A00D4B46A4ADA56858448C8246C320",
            INIT_RAM_19 => X"60AA49CA9D94E8172E463FF8D803995E9426B2A05CB2B28809F92160416ACAF4",
            INIT_RAM_1A => X"AA45A06C8D0001126D000000528080198C108493E110A000810465AC032916D8",
            INIT_RAM_1B => X"B9948B40DA70541111141494AD17555AA802D0350AADDDDD092AB46C28A454AC",
            INIT_RAM_1C => X"041554A807851E2884115700860D541556002E04020280A0B80A094B430A82A0",
            INIT_RAM_1D => X"921406200840C28290808020A053B904480A811516B5EA08F3612E80554FD851",
            INIT_RAM_1E => X"489122F4F5265C343D43B551408D777B449448BAFD005331151D85A014089242",
            INIT_RAM_1F => X"87C0BD55408F24001013BBBBDD75D75D77FFF27B5552EEBAEBAF46B555570224",
            INIT_RAM_20 => X"457084200F6AA61861804A44210840006828A281A014009120411E2228042002",
            INIT_RAM_21 => X"35D75D72AAA0090E79E789C58182208101F112409CED1640336822B820820068",
            INIT_RAM_22 => X"5C1ECD00E6AA1C44212678AEDE81BD158854210801492D044104100018888407",
            INIT_RAM_23 => X"594CBD3E06D76F052D555513AC9594B05544A0D406CAB264705097103939D72E",
            INIT_RAM_24 => X"A0944A42A4311405E3D0A214548850B1A410148501B1AD032C418250C6B94485",
            INIT_RAM_25 => X"9116C00070FC3F078F0B01040090006602030315D29546A51D4D7AE2231A3468",
            INIT_RAM_26 => X"9F255152AD6A54C929546100156A8AD090C20720013EF0B4B503731A44201448",
            INIT_RAM_27 => X"01008B00AA92124AB45B65B096EDB6C45CB311226022A2AAA902200E94A51025",
            INIT_RAM_28 => X"12A080940103101010103A1D445802400840831642200C2202002249B0241226",
            INIT_RAM_29 => X"2085458020355611E4001049208AF0450A2823A86942D2080110028858008A6E",
            INIT_RAM_2A => X"2054A32488048902240A2061232210808822F2D318E85BD0B700FAC694C0AE80",
            INIT_RAM_2B => X"800550A0014520080680106A80017000372CFBDFE4B58A4A21824438194CC130",
            INIT_RAM_2C => X"52109AC950685C2A8D0A8010909211AAFE925EA140181A042313080A02405736",
            INIT_RAM_2D => X"084490090140838202A706115A2855389A51C9A711800003541A110626582C01",
            INIT_RAM_2E => X"25184884AA01458208048FC408418C525220014B48E12AAA088095029A0AA001",
            INIT_RAM_2F => X"5A86E283EEEC38D4932A95195043C81319388B4A0D61A0A08028072A24B046C0",
            INIT_RAM_30 => X"7836CB9DF0E2E05A3DA97029242521A321489A10D29801E97A1294A52529D001",
            INIT_RAM_31 => X"D2AC5D76C3424BCC83A55880C59862215412B5C36A44004AE0A09060962A2E16",
            INIT_RAM_32 => X"D65B265CA20942094958309548AF4D34BA1815B3426804010AA90BD55A569A12",
            INIT_RAM_33 => X"5498F26721A24916452C12A8528052A555555B4DB4D481289DF90E5B495B428C",
            INIT_RAM_34 => X"4BB555261290C90A086924AA210C08A410100D14500D35D0A89281524928BFF7",
            INIT_RAM_35 => X"504041411BEA98F5F5150D24924901C8A64EEA882062022E5123EC9000429069",
            INIT_RAM_36 => X"60049A241C4045FCA4CCA3B2E449080002896A140508A6180003440C4A264EE9",
            INIT_RAM_37 => X"E4A5A4CC2D486408C9088C66367815B181F371844E90D134F15A87268D732280",
            INIT_RAM_38 => X"054C8188CD898509103C80950249EAB3A4A6ABA8AA51313A00E5E8C0A82B4868",
            INIT_RAM_39 => X"A524111485499B54044441A6F2A80A8A28098A4940020400128C539894002080",
            INIT_RAM_3A => X"8C4A6313618F04ACBC92030021C44E24CCD12D21869081C2036124FC16624849",
            INIT_RAM_3B => X"C01091B8032000024082C52235033080D8140C6AD89AC1502490515C23582C48",
            INIT_RAM_3C => X"AA423380085442071A80A2851AEF1480659BABA9693B94848017AFAF96A0A082",
            INIT_RAM_3D => X"809025248214E003244434532064B209A124B2A822844660129A26E5C9792042",
            INIT_RAM_3E => X"4812B9A66E8031014034A000006441056A09520411090031820908CAA25250A6",
            INIT_RAM_3F => X"180020507EC92530485E28421A0B4004805248208A5F52945294BBA84807A182"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"00122D200000191404BEEEEBD4AF5555DCB73ED65ABCD6BA93A56BFB4919D824",
            INIT_RAM_01 => X"110822411114482102912242088912AAAAAAAAAAAAA0AD365AAAB4AA9AFD7570",
            INIT_RAM_02 => X"8820824420422421110442224488944108922449249249249E9F891151242249",
            INIT_RAM_03 => X"5F5F5757FDF55575FF7DFF5DDFD5DFFA1084090104104408104210088A210420",
            INIT_RAM_04 => X"00800004000200040010000400100080400124DB69B75FF57DD775574775DFFD",
            INIT_RAM_05 => X"0441000100040000804000800400100010008004000200101000100200002080",
            INIT_RAM_06 => X"6809A705D1746D7A5BD6DB6B59652642C00251525D5C04000400040008002002",
            INIT_RAM_07 => X"99A2851D2AAAAAA36ADAB968A2AB4CDD7A8A1B55654495554B19308F0B1C6EE4",
            INIT_RAM_08 => X"AEEE5552A97AD52C3BA2BAAAAB57557555D926CAE4B456ACACF55552559CBCA5",
            INIT_RAM_09 => X"6A514A057766C9304C3DD5CBCF542F9F775D546202462AAAAE554AA9D5555A6E",
            INIT_RAM_0A => X"196404ABA5D5F55555D55B6EB972285B6E6B55555AAAB52AA4D4A93E2FA5AAFB",
            INIT_RAM_0B => X"A92CA5E16806906D17A745495DDFD705578F82A076570B15915698AAAD332AA7",
            INIT_RAM_0C => X"C01109585965E6DE2D54AE62E76CD821038058779CBBBBBBB3322162566E8AAA",
            INIT_RAM_0D => X"14E5DB89EF74AAAA4A8E58D6B8CC963A95558AD4555681EB5AD71CAF5254E4BC",
            INIT_RAM_0E => X"C52CAC9B66F65995562A85ABB06109DAE8151045007555D54D82173BB488F41E",
            INIT_RAM_0F => X"1A32CBB602A25555552AAB549552BBDCAAB55D95572C55896EAB531555555568",
            INIT_RAM_10 => X"66738B12AE73860EBE592574DE5EE4F681EB4B9C25AE2C8655CBED244555BB9D",
            INIT_RAM_11 => X"AA8AA8CCDB4A2A5555580059960B9CFCF822AAAB955ACD976D4EC996376CC52E",
            INIT_RAM_12 => X"74EA8656CE55654332C75C1445D000045638577C66AAAABE99155529200004CA",
            INIT_RAM_13 => X"9231560924E5086BA39576EAAA8B1646A1B222B02A055C166D155C9C8142D6B5",
            INIT_RAM_14 => X"962E759956C55D755555D872152A4CD9F3ED39CAFA5157DF7226BE6442828924",
            INIT_RAM_15 => X"2BDA06B6CDAD926E9A677712EF1738DAAAE04D0425CABB2A955DBC557559AD21",
            INIT_RAM_16 => X"942351F5575E62C42B98142C6EDA35F4C642FDD55562AB159CA82C80301D9147",
            INIT_RAM_17 => X"D55502B622A29695555556B9685555DDDD5CAAAAAEAF9DC657E2C555554AAAAB",
            INIT_RAM_18 => X"969555544B6A194A239284A90C8ED746405C32D4096A1D6AD5DD0A6A65150AA9",
            INIT_RAM_19 => X"9887A2AAAA53555556AA9D76AAB1A6A6AB1D8802BD717155936AA66B938B0AAA",
            INIT_RAM_1A => X"CD8A5313A2E6DCC492DE99F6CD5726A39996A915BCC90ED555549A531718AEA3",
            INIT_RAM_1B => X"221294A424F5AAAAAE558B2D5297555D5557230AC553333252C84A12CB098D4B",
            INIT_RAM_1C => X"95428B179A7261517155545AD4915541555A88EF7395642A1D53556A4CD16459",
            INIT_RAM_1D => X"24AB3D99B6D215550325AA8555607641352C5668A94A15B76D1C5B3650FA4726",
            INIT_RAM_1E => X"A952A522A861DAAA92AABAAE63B28CB08B90BA45F8105555555DA555617B258E",
            INIT_RAM_1F => X"2A013800516F0AAAAAE4AAAAB2CB2CB2C800552D400111451450AE8AAAAAAC54",
            INIT_RAM_20 => X"B28B5AD5568008A28A2733339CE72AACCCDB6DBE6D89BBE7CD9AE583A234A4A9",
            INIT_RAM_21 => X"EAAAAAAEB0048B4555555F629DCD177642DCB87B4092C5804295594555554A95",
            INIT_RAM_22 => X"D6561F55115553AB8B959ECD3D5C7AAA56835AD55CAA92CB32CB2C5445555206",
            INIT_RAM_23 => X"8820763B854C192081575742AA1555AAAAB15D2B1D39099C6F3C32A5D2AAB56A",
            INIT_RAM_24 => X"1D5D6EA354E502C9BB60ED1DAF35772B5682E99AA820635CA1280C0AB9473344",
            INIT_RAM_25 => X"62C567E0F038BF0F8FCFE1094AD29936652D22B5DB757557559AF84E26E5CB97",
            INIT_RAM_26 => X"2D58B42C55D58B17462A176CCB5552E323B9C8CD087802710014CAA48B1CDCB0",
            INIT_RAM_27 => X"56297B2B0CDB036CDBCF3D9D763CF3D96544AA558B1D5555566CF8B1AD6B5310",
            INIT_RAM_28 => X"5CCB36CBEDAAAED96ED9D8C11B67DB2EDB65CCF638ECDA69A452CB6021265566",
            INIT_RAM_29 => X"C415564ACA7F2F4BD9E56532C550C49755555775F15D8412AABAAAAD156A9304",
            INIT_RAM_2A => X"30339CCB958B162CDF04F8C8C0CFCB367F4F1506B596A22D445537AF15530F18",
            INIT_RAM_2B => X"62AAAC559911AAAB3215562155577F85DC520C0D41DCF104F76D9EE6072BCAF2",
            INIT_RAM_2C => X"BB9D26E157311D4AE620954A74C14BF8FEF6FEF976DEDCCB55552BB3B476DABA",
            INIT_RAM_2D => X"D6B143D2458F1DE54AABCD5552AA955E450AAA9CAA555557E3A66AAAAA572BB0",
            INIT_RAM_2E => X"07E2EAC0E891D666A166ABD4A516B4AA53A58ABB1B1ED5B556681C4FB5541936",
            INIT_RAM_2F => X"D29CEACAEEECAF9ED88A22C3469BA9673E3EAD5B616AB2BD02373BACB6B34932",
            INIT_RAM_30 => X"ECDCEB49D8EAD75B45EFBCE9B635B5B3D9CFA61E8AF6D9AD6B1ADCE635ADDECD",
            INIT_RAM_31 => X"E3B46F76E64B734795B95A9AD5A959BDD6AC39AB6248A57318B893B9142B4E45",
            INIT_RAM_32 => X"D79AC76AFDAD8CAD919EDCF64E2F71A4D79235AC738F17912EB9E5556358E312",
            INIT_RAM_33 => X"8B22AAA8956986356B8BB2856B646B455555536D36B6D1AB1DDE2B1A49736B36",
            INIT_RAM_34 => X"A69C8DAF67D1DE2FB38DB6FAB5B33B054555315554E750DE3CF236A371B25DD5",
            INIT_RAM_35 => X"DD1555525BEA26F5746443D75D75E3B3058EE8ACB2AB5BC505101928C58E2616",
            INIT_RAM_36 => X"0C56DBC8A2ACD27B1550D5555528A59379D95E8BB1AE08B1AD7399318C759EEE",
            INIT_RAM_37 => X"B275BBA8A4AE57173A662F6E637AED7795D733957ED74B70EAA9AAD8AD745916",
            INIT_RAM_38 => X"585CE662E99CB57DC0859FA57EAC8C2DA796AAAF9576BD8A4801E452571F256E",
            INIT_RAM_39 => X"72B99C5CD7627B5579555D2E49AB4AAAAABB9ADB5FB6B1BDB6BCD7B9B5FAAAA5",
            INIT_RAM_3A => X"2E6F6738AE50AAA8C15D8A535528017436DBAE31A6DAFD56BA44DE7896E36E92",
            INIT_RAM_3B => X"92D8F7BAEF4DBB6E2B1ACD6E752A793BC2A6AE6BDB3A9B5AB6DA9A7DB77A2B2E",
            INIT_RAM_3C => X"6B6C5BBBC971466F00D53B29ADD637F735D9103BAB1BB5A91B000000C33AEAE3",
            INIT_RAM_3D => X"B6DAB5B49335EC222554A55B2264F34DB5B6E3AD4AD717655CCACEEAC979256E",
            INIT_RAM_3E => X"491B63B76CFD635A09D4E4C09BC96DB7FEAD9BB6DBB73573980DED32CB5B59AE",
            INIT_RAM_3F => X"D800D97CCEDB5FBD34008A7392AA5C1A079B6DB6DADC8B5ABB5AFB6D4886B9FB"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_basic
