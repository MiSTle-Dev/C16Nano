--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10.03 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Thu May 15 13:07:37 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_funcl is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_funcl;

architecture Behavioral of Gowin_pROM_funcl is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"FAFBD0049CCC831FDBD0072434F61A9791D00E481F1D7F81DBF61CBCC7997E80",
            INIT_RAM_01 => X"DAA10840DC0582308F5CEDDB76BDD5FBBF4790080074BA0A0601AD3B5E0814EB",
            INIT_RAM_02 => X"486D24080D34A1120ED1403D5D49120B77A664CCCC444CCCE4C343FD6AC620E3",
            INIT_RAM_03 => X"D489011E482D249A5136C341A60A0492C92C12D80C92926924C004A498488054",
            INIT_RAM_04 => X"D90CBB416CB4934E20BFEA4BFE75511FCED09E2DBB5B6F2429857C4405954153",
            INIT_RAM_05 => X"C2450C4B93862549CA248A700A8B1862108A2913243F0BDCAD3113530A215A14",
            INIT_RAM_06 => X"FC19A36F8F294F3488D59811F1CB4B0526B752714B78D2694E159A4B29896248",
            INIT_RAM_07 => X"42821F49A6987058FA07FFFD5C028A0AA2A5F7D705C299462143E529E68D6C68",
            INIT_RAM_08 => X"C7D4DF7FF47D0A52909B20A54B25C9A9E99AB00496D60A7400C5451250B0250D",
            INIT_RAM_09 => X"016041A00492D958375316571412CAE2D0E9322AD5EB7242574C75FF6A474E4F",
            INIT_RAM_0A => X"FE662D5E5DAC06D327940F65EE702982E4050415DF47AAF1829624A7DFE854DD",
            INIT_RAM_0B => X"9A94DA52388423C0B8840405C081953EDCAD4D11058755378913E35809068E42",
            INIT_RAM_0C => X"0024F0A1ADC5A3FB5FAE5F2ACB4463262049374331C26CB4B452AB43B09B84D4",
            INIT_RAM_0D => X"E5A48CE9B9590912D8D89C8020A5DD9670E228134D34FAF54943628B0E646DB8",
            INIT_RAM_0E => X"E1C6D0094E3836276871F0480565458217233087CA250EC8995F1328117934EB",
            INIT_RAM_0F => X"A898596E5D640A000A79402C0108A53C1666932E932E834753BDE7E3CD027662",
            INIT_RAM_10 => X"BA33ABA0D96AF4BC1F3F317858696FD48B69A25B4D908D7517E1346A7C0DDF14",
            INIT_RAM_11 => X"AD80C82D5100919724059439400D44A22A12455AE0A1005FA2ACAA6A741D1084",
            INIT_RAM_12 => X"AD6B7B50ADE09389147282F68D9EF6EBA7245214876DFA051EA5F439EF2E6F22",
            INIT_RAM_13 => X"6D4E855A0DD40B705CA20B2876A90165264100D921900202654094806486558F",
            INIT_RAM_14 => X"42AF329A498232AA2E6100B5644425017A410C86D105A616E95955197378B340",
            INIT_RAM_15 => X"92A95400A28A10A002208CFA82D29F55EBFBDABA432D32946762C02510581258",
            INIT_RAM_16 => X"91F2D3DD9B49049B42A2A65795852008214005228493124014453C9681640802",
            INIT_RAM_17 => X"084501500894008B68D0A8BB044A052E3CB2505C9185D3D4AD161E0D0A050D4C",
            INIT_RAM_18 => X"A91EE1EFA99538104029A944E050A402783428A9EE010687B420F50F72534169",
            INIT_RAM_19 => X"B252461726280D1001A00229AA6094B26281A3540D404B431609CAAD23D83D4C",
            INIT_RAM_1A => X"1615802F2E20FAA32A8AD02462D10493469AA86806AC54926869143400A2D528",
            INIT_RAM_1B => X"9994402688A130FDB5FA240E18B474DC8705009406E99C6801A808A204189400",
            INIT_RAM_1C => X"13497915212EE68EBD1A37FEDBDD098B5CA22BABBA16C55C062C6C7E2A5DAACB",
            INIT_RAM_1D => X"74213291BC92273B0D1C839D51B128D8E09B6B8665D6B8D5C6BDB36B82185653",
            INIT_RAM_1E => X"D8EC9F63A840CA68AB16EA402582D5815ED4B49A5934B99A45A31412E66385AE",
            INIT_RAM_1F => X"8D31B08E98A636DB6DA2C116ED5EEBBBDFBB2F1D75ECCC7DFA6484832A64EC9E",
            INIT_RAM_20 => X"F9C6FEC412D825BC6BEA6BE565A77EF35F35F2FB4C231845BE8DA3FAF6356306",
            INIT_RAM_21 => X"4009EFF589BC6D9B4490682051203F51FDE7D4C975510556FDED38956AFA4AFD",
            INIT_RAM_22 => X"7E6D95E2BA5D55A900ED78205356F5665FDFEFDB2F6FF7EDAAF5571AB8090482",
            INIT_RAM_23 => X"2A052D90F6FF6F608B5ECCBC38C920131C09AD7A3EE8DFB9B6BFF271D52402F0",
            INIT_RAM_24 => X"01E610760157515F078D7FA29CDE4F14E526AC3C4445BF8CEA2BC3AE34015BE5",
            INIT_RAM_25 => X"BEAF6DEDB96B7EC8A3E046D36B8649459B0D61AAE85A486AD7772BE1CC6A60E1",
            INIT_RAM_26 => X"E1684EC1301247EEEEFEEBDEF4167EF6EE020D726B80BFFDB1339EF5153F9BFF",
            INIT_RAM_27 => X"E55F5ED789A8D89CFA9AB7A4ED5DD99BDAF37D77EDFF57CC24E21556AAFBABFF",
            INIT_RAM_28 => X"30DFDEAAA0B92497D20330C49885573716B5AE3E26B7276DAFC559996D7B9DE4",
            INIT_RAM_29 => X"105A040441410543430FD08BEE53E1CF15A4796A1237774FF5B415D3C6FEFEA1",
            INIT_RAM_2A => X"609D1FA5D28B4B791EFBCA23720446E424119DD4989A982132024592582EDFED",
            INIT_RAM_2B => X"4DB40A502E823556A836A4A54388925A23275688ADB60A5604BEA1CEF7A98ED0",
            INIT_RAM_2C => X"520A7001F8338C3001F8B47068F1D9F2CE8E0AC849DEEAFA1A4A9449465232B2",
            INIT_RAM_2D => X"93D6ADF4A7E6B6D6FD496E65FEF06BF6555B59435C611AA543108B63A06AB491",
            INIT_RAM_2E => X"6ECF8151060B867A05C33D059626EF238219135A956A2BDBCF76B76852EBDB57",
            INIT_RAM_2F => X"8913A0BD7FA7DD4D4B7FB513BC9040F202576AAAA92922A124852023E48095DA",
            INIT_RAM_30 => X"5BFFB34D7FA5377E545A84986417BE72ED7B2C39ADD665F524CAC9A447DD8BE0",
            INIT_RAM_31 => X"0224350870456011624885605586BFBEAFD7CA23D6F5EBF9F655514AC4EB5FD3",
            INIT_RAM_32 => X"ABFE511F991D995EC0475F76611F9287FA606E2384A96310AA589D087E514017",
            INIT_RAM_33 => X"DF6C20940275E37A04240E8886E3ABA001011875FB5B819C20153023198056AA",
            INIT_RAM_34 => X"D55DE746657BBCD4B78AF15E1E964AE532011101119DEF31B6FB17FAB3BDE746",
            INIT_RAM_35 => X"E98F55E8FC9B3DFFF564FEDA1D79F84BAA91925D50A91F1F7CD4ADBDA7BFB421",
            INIT_RAM_36 => X"61ABF8AFEDFCBDB4EB750CC5E204D9BF8265F4D94413B650646886BBB934434C",
            INIT_RAM_37 => X"3EAE78EBC3FA18386386B8019754F9BF57EAAA54E9E8F0C70C70D7100F0D3C82",
            INIT_RAM_38 => X"70586364AE5AD824D5CB5B448FB7ED0424762F3AF3B5FD7EEDF6EE5F647423D5",
            INIT_RAM_39 => X"CA93F486D82E6960A696ED76AFCD849A1829A53D7FBB6D57FB77F30CBEC06869",
            INIT_RAM_3A => X"22FCDDDDDDDDDDDAB17E4D3BE45F91D7533AFAEAFAEAFAEB5DAC75AC7E5515EB",
            INIT_RAM_3B => X"9AEAAE3AAB83F5FC5AEA81797F276F37AC2E680C35C3D223C0C35FB7FAFDAAEB",
            INIT_RAM_3C => X"0FC13C0E053C7E8E9C93F53AC28E9A43FB68280BFDA0A8F7FBC5B7FD7B2BFD70",
            INIT_RAM_3D => X"C91FDD417A92F5042F9F1F3E4D3D59F74CA002478BAA5F27E9B7AACFBA650412",
            INIT_RAM_3E => X"3C32C1ADD3931AAC5635D71C5CBAC1DA97D22F56B881648FEEA25EA4BD416143",
            INIT_RAM_3F => X"031C32B7D7BE56081C7AD3AAB48BFAA9DF55F5BD0EBD57F5FE9B64C164B05216"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"002D6FEEC600D074010242429C404C0154A400120240DA0501014588410A9580",
            INIT_RAM_01 => X"88AC8C2BAC052282804468C65024A02904092828141017FF0200C68023B64894",
            INIT_RAM_02 => X"0001A65118841000A504A8890A0000A400A02AA822AA2A2A0A82200A85284508",
            INIT_RAM_03 => X"62024004114926500D904B4080820004DA4082D26812924D24DA6D300B01B040",
            INIT_RAM_04 => X"CF504941596B6C8400ABEFB4EE2E77FC030209D6A9AC178C86A5162C646F24A1",
            INIT_RAM_05 => X"23860290E04148B02149B16A9015490094A2A997BE66ACA85270845A112DA804",
            INIT_RAM_06 => X"EE3A210A56002210CC811533E2AE4A802C5222E846703A662D1A4092C85A9488",
            INIT_RAM_07 => X"C481636084D1B19B1B720A2282820A2A2A85DFD7918A29956804C004421638E9",
            INIT_RAM_08 => X"880001221D08C2A0AA2135288140430302C12C696912562C00804026102C4108",
            INIT_RAM_09 => X"404201611269361100000989004520098211108002841180902252C634008018",
            INIT_RAM_0A => X"08B064018A44A98D5C6150284413412C0150DD60452046082828901148402500",
            INIT_RAM_0B => X"21422003AC114910114C6A00418FDC294219DE30C165081032106948832585C2",
            INIT_RAM_0C => X"0220A8C10943224912961A344340A1AB0302C00844A084401614142815511900",
            INIT_RAM_0D => X"140A112244800A502082891ACA2882014441811411490000000252860B204128",
            INIT_RAM_0E => X"22700A04108982490E9058A19240408225225004800C84986028000100844200",
            INIT_RAM_0F => X"190022143606C0084C304220001046191002180218020A028CA049046011A300",
            INIT_RAM_10 => X"162083199BB1206805111C963512C214034C80D16522080D094DD9B01406884B",
            INIT_RAM_11 => X"40028040D4282FA1042181128400022100892210CA0D12C308840290014B4834",
            INIT_RAM_12 => X"41CE10224124890A20841028502014490200218020143091D419209053111411",
            INIT_RAM_13 => X"42080281290C103584014302241108600C821001012208C80808040049840102",
            INIT_RAM_14 => X"4404228A2092411080D0C50041800A28C0092902006D32430F8202D888A44201",
            INIT_RAM_15 => X"9420C44060961061100893110D0908849000851042517FE97846000910909212",
            INIT_RAM_16 => X"000408100630C0000060652C6228008602228800814422842A86198022232ED5",
            INIT_RAM_17 => X"030000369101CC45021442492D20B0B0A002850401205A8105028840A080D010",
            INIT_RAM_18 => X"C04B694104F810DA04030480960C0AC82D0282114400C5A0233B884A28B2C258",
            INIT_RAM_19 => X"40000481180A0B03416A22C30230A01180A162040B51CAC0632A9040016D0827",
            INIT_RAM_1A => X"40A05A0152400004844102C10000410C441008442421882188402420130C8102",
            INIT_RAM_1B => X"0D3298A4016148002290150590C4A4F63021600C22A0202E056C2010F28121CC",
            INIT_RAM_1C => X"1F00494DCD4210C218D0800A659274A40140D4A4B41AC91B5850A0B6422A85A4",
            INIT_RAM_1D => X"2B952116A480101A2049892001230090061240A0310100C804890600A6C10500",
            INIT_RAM_1E => X"41240402092AC0C8011C1088210002108000432180350A40002D18D4210C5810",
            INIT_RAM_1F => X"858C24D4892812492483113024045009000020202048622A00C802190AA42512",
            INIT_RAM_20 => X"0D1900684DA09369B4813692531291A936DA4C180D3582AA8184192408108102",
            INIT_RAM_21 => X"509920A050880100250080040204A006281889A4C0D6D8282A58826A00115200",
            INIT_RAM_22 => X"FF289202404218C3A2C10ED982A3583F204180841020C04210082019009A60A0",
            INIT_RAM_23 => X"90A49888CB08226028251605102030C1C9040014838089001B149B50089C06F7",
            INIT_RAM_24 => X"4042010998A820500005944C5AB0C762D7CC4D2101402080CC32433620926049",
            INIT_RAM_25 => X"100082405600200810190085008F6882010A60738431901CA46A9A604AC54002",
            INIT_RAM_26 => X"04C0B579C060285005002D2260820401421A2D134A0C008B18A8D09000C24404",
            INIT_RAM_27 => X"738F6F308BDCAD18FE28BBCC3539B6DDBD7A7FA7BDA7991794E313FC05015400",
            INIT_RAM_28 => X"305004010C053482CA60C0130A05A03171DDBF6B37E2BF1C8F2B693BB11974E4",
            INIT_RAM_29 => X"29604A200A0A2A080820D0C04210018DC5B744224834200080008512A41A6445",
            INIT_RAM_2A => X"6C0091329006A0D46090900C24D12AA8067428A9550F1B00360020860B098492",
            INIT_RAM_2B => X"49A602040048508A8A0100509104C106186A410604484A820900000000020404",
            INIT_RAM_2C => X"19B3B2C84CA516B2C84C249ACC129824C4940D630090505021902512CAA4212B",
            INIT_RAM_2D => X"4021025000220900009F76652103452110202258030D401A310042E5A0442680",
            INIT_RAM_2E => X"40000CC0180A4024052110000002002181843204095008201001012100000409",
            INIT_RAM_2F => X"851590AC85280123250600D1B44E3ACA162208210565400C307481659085C8DB",
            INIT_RAM_30 => X"801245969000222481081200652550441014B823148A6520E0D21502328A6229",
            INIT_RAM_31 => X"108D3661A12A138081C25A0249120A1B01836D3800D9832DBE00221001000485",
            INIT_RAM_32 => X"4A50908A408A40242C220A2100892E425B53082D052002010258880025054402",
            INIT_RAM_33 => X"38600908861898096DA2440DC0008319120328189942100DB60D1A3602182640",
            INIT_RAM_34 => X"C208B21320201108C30C61AC030650291411B211B1284A000CC01165958D6300",
            INIT_RAM_35 => X"09ED048284A061ACB4A5D6FD2A22810901044D480429D5D58A840618F212090A",
            INIT_RAM_36 => X"2CA1A45006500100002104C0002000408152A84269133798100A00028A000010",
            INIT_RAM_37 => X"250450B530A4288822801685016290502040102041485141045002C0051A0849",
            INIT_RAM_38 => X"8C0081BC0600D2A480C01A14835096D3AB22150C441A84B000A0462B42084418",
            INIT_RAM_39 => X"030420401121494594969036842116D211652412252080010101436016CAC15D",
            INIT_RAM_3A => X"35048080808888991A82099086A08082141202120202121144472447240F1521",
            INIT_RAM_3B => X"9040041001180A4400482D0C94B281A004011A28942092080429361945004555",
            INIT_RAM_3C => X"436548211816A54509D4B590CC0CDB7120010CC4800406412432012724E09220",
            INIT_RAM_3D => X"49A82924525824902306460C6D19198663740D96C00120E91A0808CC331BA0ED",
            INIT_RAM_3E => X"14141058961842420800890408002808000F0504A230A4D40490149609244424",
            INIT_RAM_3F => X"211412130695299EC84100002D10805884825059021A280050D8414A0904C4C2"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"52BF7004B40C932B8D2307027CD13E5345C68C482F451D4AFA52499682D1424B",
            INIT_RAM_01 => X"C294260FBC1981706BD9F4D7743F81FE0F4285005469AA0A0004E71A3514404A",
            INIT_RAM_02 => X"0943A4008CD806A88681422D0DA2A88A44CA802288A0A020001237ED224261C2",
            INIT_RAM_03 => X"71F1658BFDD6592E9F5B6F90DF37F27D65B25BFBF2FF6DB6C92D92DD27934860",
            INIT_RAM_04 => X"755516D034DB6D0A10705AFEA3343C30FC4061797C0305A0CF4863BB1280399B",
            INIT_RAM_05 => X"A98FBA7D635D3EB1AD3FEE113FFCEF2895A02B26AF9D4172BEEDE1BA2D7DA6B0",
            INIT_RAM_06 => X"9458CD717895A5A1E13E5FB50ADE7934ECA64952FE455B3DC255DC7EC75973E3",
            INIT_RAM_07 => X"5EA1536A3481F5569B5DF57D75755FF5FF7A0820EA33DF7F2D2D12B4B42AF94C",
            INIT_RAM_08 => X"A144035668346C5B1AB820F4CF6D0F8F854C942B694548500D0040364851E494",
            INIT_RAM_09 => X"58825A013FDB7FC89172635B73836A2BC2A984AFF1A503F2D503AD294931239D",
            INIT_RAM_0A => X"BEF28F7BDFE61BDE7EF51FAEEE4A09AB15177D5C2E32C6580BE8B5B79DEA5DC4",
            INIT_RAM_0B => X"A9FC3B4B38F63EC5E9C02E2D00075656B4AF575B4CA34DA51124D2D418020A02",
            INIT_RAM_0C => X"12872B62165800B2CD68050AAC526946816BD22A5F4AE076B473F62B00CEB3C6",
            INIT_RAM_0D => X"508B5D4BD1EB61E63847147FEBEDE7B250D0EB0514DD7BF76944A5B01604854B",
            INIT_RAM_0E => X"8AE6A31516A137677E74F068D565E4326924D2E9AE39CF08FEF7956BB3EF7FA8",
            INIT_RAM_0F => X"F7A951ECEF6C8C6B4EB99A84021D675D4200B220B230B3675FF5E7B2C563F227",
            INIT_RAM_10 => X"3831EA91B6D2D5D8BB296D6CE969AD06BA682E98417E8BCD16CBE97AEC5F9456",
            INIT_RAM_11 => X"E512466527245FDC6DADBF68DFC5779000692DCAABFD97F6A33CE27ED4181CF6",
            INIT_RAM_12 => X"E2E72F70FC98BFC11042E7FE1C3DC3A38D6CC11CADFF6ABD9FBDF43BE6EBFB56",
            INIT_RAM_13 => X"235E2DCB25CB997F71B75B7ED19B6B6F7A337C5272705E8AE741DDCC9C52D58D",
            INIT_RAM_14 => X"2E0BE1043C22E6E2BAE8DBD341EE1F8BFAEE25669709A01FAFCFD5D75FD5AB49",
            INIT_RAM_15 => X"2040168002C020022812DFAAEFF3B5557EDBCE2925C039E17726F118C9A84A28",
            INIT_RAM_16 => X"D32753D50F795EB2C270F3DAD6B1F08AF08AA03243B7F0D768275D6286222468",
            INIT_RAM_17 => X"6E5551379F9FDC1A60D0A2A0296EB7383D327FD0C7AD13C0B1188FEC2FADD40D",
            INIT_RAM_18 => X"E157EDE6EFFC1B9F613F9D80C4D8FA983FB0BFB1E6B04623F211554F3B030EE0",
            INIT_RAM_19 => X"F6DA1EB47723941F728280BF8CE11687623A851D9454A30E5E3176652AF9B5FF",
            INIT_RAM_1A => X"C69D7A390804EF9DE6214FE1EE57673B2A28C4A59E197CE764A1E250CEFEC67A",
            INIT_RAM_1B => X"FC1248360481BC4C77E1AA68A055F16CFFAC36002E891CEEB50E2AC0728F9FDC",
            INIT_RAM_1C => X"8B5D5254A41C2485A492B5BD9E442DAB54A0AA3A2B0845D554A8786A2019A3C2",
            INIT_RAM_1D => X"7515B0951541157061508A144A03242032F95982DD52EE57710C8D1981494341",
            INIT_RAM_1E => X"807805429F3ADFA19B1E8FDD820A3DA16A59DEAF7B907092EC8A0851C24A143A",
            INIT_RAM_1F => X"0522858E0D44124924A110962DCB2392FE394FAD21654A7292C005CA54897807",
            INIT_RAM_20 => X"481D5E48DFF9BFDBDF79CD3EBE94EDEE6BAEBE99CD63082125048BDA54156142",
            INIT_RAM_21 => X"8005FF50100C2509338038A8140B37374ADFC17FB4859C6E7394F3FBA0F51854",
            INIT_RAM_22 => X"1C861F1AE15F1CEA80A9D4510113DD577E734AD6FF3BAD2938FCDDCAEE292F03",
            INIT_RAM_23 => X"3997F41C24924B72AF4F5F9C307884F39D0D8F29FD7F7384FFAFE051A0B407E0",
            INIT_RAM_24 => X"40B41B5F8CF51343634DDF6B849EDD5C252D29F24D04B94C6619C19DB6617604",
            INIT_RAM_25 => X"28AF6FE7A72DCF7BB751035B62CD4AA1C02841D222B5707561192FC1A8D890F1",
            INIT_RAM_26 => X"2A00445714501E2EFABA3B56FC107F9FA3D8447843C5DDFE9408A7FCB6FEFFDE",
            INIT_RAM_27 => X"B9AA677DFECA8BD9E7DF68D7A9B93BF0D4625F7CCFBBDC9401A3AC0001414155",
            INIT_RAM_28 => X"925EDE2AD435BE87EB61F8E78B42F3B2BAF76BA3BF67FD2ECFDBFBEDB53EBDFC",
            INIT_RAM_29 => X"39385904626007606007A0F9A259318DC1FF3619603B7F0F47D62419A0F7FA41",
            INIT_RAM_2A => X"5D94D947A09AC3583B78DC45D295C0A80767ACF1D11D1569A8D314534F6B4249",
            INIT_RAM_2B => X"430E00006659B444AB04F025434391142B84858A2F6F127604AA8944B5294F50",
            INIT_RAM_2C => X"0B894A22FE039E0A22FE047A1C7B30E6999EBECFCDFE59C88E7E1404A6893BF1",
            INIT_RAM_2D => X"8AF32EF2A568BED2D2BD388D5298EFC2876060FE73CC7E3F70400163102E0E41",
            INIT_RAM_2E => X"5E6E1144A3FAB74C7D5AA6048F1CE98723EF295E73533EFBDD32F6DD728B4D5B",
            INIT_RAM_2F => X"4A3069A34A62D2FE0EF9B4C302B7DA16155173EA4A6A42EFB5B561522D0554F3",
            INIT_RAM_30 => X"DB7FB7DF7DA5277E518658065CC33654E72C0A2B29908D5166B851B45516A2FF",
            INIT_RAM_31 => X"54C233E8F5974121E3D32F214C1955BF8B974E3AD0FDAB79FE1D4042A0AB4FD7",
            INIT_RAM_32 => X"BAA28152A150A1CA0054904AA55794A796089B0F673CE2042A7898046E5D8057",
            INIT_RAM_33 => X"F3AE0484853DED4760254A855231EA910902903DF508D4ABB090281548DF50B8",
            INIT_RAM_34 => X"4208A0122703801CE38E71CE0F81C228D400A900A894A575FA9F9FDF9A94AD57",
            INIT_RAM_35 => X"53CF5FEF690B551DFEBFCFFD9C7BE83F05A6FFB8252C9292D606A7BC65FE9F1A",
            INIT_RAM_36 => X"EFBF5CAD6FFD9494B95828A5F060DFEFAD216413DF1409F57C50A5A0A22C52C0",
            INIT_RAM_37 => X"BA9A287BEF5A30B0C103AC1D807CEBEF7FAE2850A1C0A0821820759ECA047692",
            INIT_RAM_38 => X"7E48076D000A1024E001424486BFFFC7A65C2A1EF79FFF6A1866B8544CFE625F",
            INIT_RAM_39 => X"D1A2D080550550559507FF073E455694154541ED5A1F7F3EFF7EE3A43EE27051",
            INIT_RAM_3A => X"E6EEBCBCBCB4B4BA93776B2944DDD945115BA3B3B3B3A3A10C9B529B540E39DC",
            INIT_RAM_3B => X"0EEAAE3AAB8795EE7A52A471EFB5EF2FE038650A90A1A021002F6FF6DEF4A6FF",
            INIT_RAM_3C => X"F67A1C0510387E2E1C21D0380808E42BFF6821AFEDA0B8F6FB47B7FE5BCBFF02",
            INIT_RAM_3D => X"AD3FFA0D740AE835C70E0E1C7A5D1D047F5ECB04EA295B43D0B688E823FAF24A",
            INIT_RAM_3E => X"3826ABBCE7D75CBE161D573C940A3DF08145BA153AB9D69FED025D02BA0D5577",
            INIT_RAM_3F => X"2608239ED5BB75144428D2E39D89DAF9CFE7FCF427B7D6B7EFDBC0EA7DBC84F4"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"E71BDFFDBC71831CF6C41964592E2CACC0D83240D38DBE8F1294159282520A49",
            INIT_RAM_01 => X"1A89084AED987BA80650198E073FECEFB7B9EA204759B7FF0205AD0D1A28A89C",
            INIT_RAM_02 => X"6806A6A9E6C8CFFB0353806706EFFB1C66C46CC6EC46E44644E5B1066CE6DF6B",
            INIT_RAM_03 => X"05ADF7833CF24BEDD3FFFEB0EBE5B24B76DA59FBD36FFEDB7DB6DF4F2592DEBC",
            INIT_RAM_04 => X"755DD6F1471B6DA0110EB4EF498E3110CCE0C35157E2CD801100205243105C81",
            INIT_RAM_05 => X"4D929416694A0B34A60B600311104D0A152A222EFACC7022136CE0BB364CC6B0",
            INIT_RAM_06 => X"84104E45DD00C4A0E03CC7B1531F5C516E0308425F68527C00515214C28850A1",
            INIT_RAM_07 => X"80B2366FB48DE4CDB32200AA80AA28022AA22222775AF9612045A0189403FC48",
            INIT_RAM_08 => X"4698CD5BA9D5FC3F0B3B0071542ADEBEAC97618B6B6780F02245190007180066",
            INIT_RAM_09 => X"0624048202FFEF22E68C45EE65D16CEF5BC524F454EF71C41E44CE718DA6B556",
            INIT_RAM_0A => X"BEFA8F4BFF8B35EE7F7A1DE35538252CD816A169F4450AA58B56B7179EE62DD9",
            INIT_RAM_0B => X"2BE07F9A21EF144059C00FCAD80379E739C4F7EF9FCFD1B308A73F9FBC6E3F00",
            INIT_RAM_0C => X"22EA7B6CB4C1A2DB56B416ADFE341E4080F3D46F5A2CEDFF30F1144EB045ABFF",
            INIT_RAM_0D => X"A52F77EAF03680B17F4DA4DF83E15BED75E26E571DF9EEDDF259B58354652998",
            INIT_RAM_0E => X"62C6385F16B8350A78A541AB1653C98092092072E618F6486FB19F4E22B55AC3",
            INIT_RAM_0F => X"DE3152AFADB8DC589E7F86E08994CF3F7024E04EE05EFA028FE8FBC501F1E404",
            INIT_RAM_10 => X"9822F7A2FEFBF95D2FBB79FAAD7EB754F301BCC30DFD2E919FEB7D6CBE95DD96",
            INIT_RAM_11 => X"08005C0865489FEB4C220A8B1508730E4C482A35F2D1A57BC33EE8B9890C4EF6",
            INIT_RAM_12 => X"732879BA677CAA780819757FDD3B316BFB59922B48BFBD29151D72BEFBD17DC5",
            INIT_RAM_13 => X"2C7A8A10057B023DAD3144151723088292E014821C939555AA9C6C6324A5AA37",
            INIT_RAM_14 => X"528BE71C1DB2A44CB1A0014641C3C692BBE604C09E2C060EEB56ED1E8BE14840",
            INIT_RAM_15 => X"14A1160488D010800C22D6D50B43CAA17C52D6AA59367EE15DC0A02716481449",
            INIT_RAM_16 => X"CA61829C37BE1228855555EF7BDA933092C0B91038CF02059CCF3F542944489C",
            INIT_RAM_17 => X"111862414E2A10D568C142DB397CFE2CADC2AAAD694ACA105CAE11A1BD4A1507",
            INIT_RAM_18 => X"AE5E844955B554450555374832A554504686F548510E1C042522AA82808610C3",
            INIT_RAM_19 => X"F9BCA52B5442E47D5C8286B53C870F35542C897C6454B81158707C8853D48AAD",
            INIT_RAM_1A => X"862AA1533659B6D7E8B3EB81FCDE0E2A134BC335014565C54337C19882D29E12",
            INIT_RAM_1B => X"EDA090B48400DC1C628B0C530815B336ABCB4190486A2DAA098A436284562A10",
            INIT_RAM_1C => X"867D7A5C0C366408C51D56BC9E67552D7758B0383800DBFE5490383E0C4CE9E8",
            INIT_RAM_1D => X"7001A4150542355B655DAB8114F00BC876F17212BDE4D486A538B93211C94153",
            INIT_RAM_1E => X"CCDCCFCBBE5205233054351064906AE95BD45AA96FA0D993E90B02C3664AD539",
            INIT_RAM_1F => X"8536B58419C21249248051B48852CBB1DEBBCFAF65C4CE56B3C019DB7468DCCD",
            INIT_RAM_20 => X"38DC2ECFFF7FFEFFCF23CF37B6B5E35E7BEFBE32A9611044900423DAD0152102",
            INIT_RAM_21 => X"490569449938D3269615A93A1C0FA867BB3C916DA583DD1FD6B5AFD4C8FE4229",
            INIT_RAM_22 => X"7FAE8D58A90555BB10F5E8A2A2E6F76FDAF7DC626D79E63128B49A90D4F86293",
            INIT_RAM_23 => X"2A17B5452CB2C99F0ED2960158B090239F440B5A142B0FC917C5E830880005F5",
            INIT_RAM_24 => X"0094033FC47064054489CF2800DA4540050E0845100B6AC1775DC5DBB06972A0",
            INIT_RAM_25 => X"EBBBFDEDAF6B5B90D1A2A463CB8DE105B29541DA68B91877390C0BC194E220E8",
            INIT_RAM_26 => X"AEFBAD5ABFDA5AD11004DFC3D0B45A368B410410028440B6B531A9FD37F576DA",
            INIT_RAM_27 => X"318A77719DFD5C72630C2CA5A15D31F1F6E74DB6CD332B305A5F0547855403BE",
            INIT_RAM_28 => X"0696DE83140D0C973A03FBF7198577B3B2B766666A2A2528AF077B3FFFA81EB5",
            INIT_RAM_29 => X"42008748F9F980B9B9806420ACD042D6F4DB0B60B20D4D6BD77201CAF0AD9EE9",
            INIT_RAM_2A => X"B015024523118E31EDB9B5DDEEF4CECB3553A9A7191E8D001A401861940F56DB",
            INIT_RAM_2B => X"4FBE4C774A951D12EE261097178F831E3BC2870EEB6F44B6B9BEFF6FB7E94ADE",
            INIT_RAM_2C => X"12802849B4310A3849B4362878D2F1A49796BCEA85BCB7221BDAA556C2AD2B7A",
            INIT_RAM_2D => X"D3D7FFA4F3E4F7F7F457B2CD9CB2C514C77171F776E85EADD35CC8C1B44ABE91",
            INIT_RAM_2E => X"1ACA9506A9BB279E5D93CF09172CB325ABBF1A5EBF7A5FFFD5E6D7F873AFDFFE",
            INIT_RAM_2F => X"4F3349BA52E6F6FE0E79BD858EB7D236235673EACA6A62EB35A562206D0895BB",
            INIT_RAM_30 => X"FFEDFEFBEFF077DE74D82C8C38D5C87C394E0E7B80C2CD9674780D80196723DB",
            INIT_RAM_31 => X"1065A5E270CFB805E381874041CE0AEDAAF5E79AD66CFDDCDE1D5D8CB4AFDB7E",
            INIT_RAM_32 => X"3B2A9065206520728019E59CA065843B2E21BE0EC7BC4199A872BF087F9D8587",
            INIT_RAM_33 => X"F7AE24208B5EEC3D4C2814821042F7A24845005EED01101730A0520941161C33",
            INIT_RAM_34 => X"00000000054EA775E7DF7BEF67DDCCA8D460506058842115FABF9EFB28842157",
            INIT_RAM_35 => X"F2C653E9A91B6267DBDB312C3FFBEC0FB083FFDD80251D5D58C2ABEDA3B7B56B",
            INIT_RAM_36 => X"8E2944631D345E5CE3C608781AA40EB5BA14309BDE1CC9F616F0EF3B1B78779C",
            INIT_RAM_37 => X"B82080BDD9CEC101040442401272E0E7738BFBD7AE31E2082080885CB601DC40",
            INIT_RAM_38 => X"4383B16B2A9F40122553E8024294A5000170782F7834A5282100E2F10003209C",
            INIT_RAM_39 => X"6CDED4528622101921033F43388866C4864841D9B6C7EBEED70E98A83A3823F9",
            INIT_RAM_3A => X"700435353735352AB802022B760081554227AFAFAFAFAFA8011A561A54AA294E",
            INIT_RAM_3B => X"44FABF3EAFD6B4E47E93CC51E935298DED3B144300422040688BEDFFFE704D45",
            INIT_RAM_3C => X"A0BA7D40C5FCFFCFFCA7F13882F3761AFBEA486BEFA92EB6FB75B7FA5B4BED46",
            INIT_RAM_3D => X"0988A26244C4898961E383C7B62D0E59BE48B2796EBA7FCFF3FFA872CDF24193",
            INIT_RAM_3E => X"482062F5258714F416221F2C6C9A85409350A8112C8004C44134913122621904",
            INIT_RAM_3F => X"802022B6FDAC5A28A0537D0D49834FB15B5DB5B60AD4B18C25D2C06A5DACD4EC"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"A528401DC6B6CB04635DC1249E264F84DAEB86C9D2271A8D2420102D45ABFC00",
            INIT_RAM_01 => X"0540511089320C0D1026008309249688043513452064D10019509454AA69BC94",
            INIT_RAM_02 => X"08E8A603013222205C38351BB882204199999191BBBBB999B308401800108010",
            INIT_RAM_03 => X"A4D24918926412596D020900B08B6D261B4880906524DB4D26DA6912D301B147",
            INIT_RAM_04 => X"D23372435D7924C800AAEFBBFB0A56DF3FFF155A28920D08487B800488436372",
            INIT_RAM_05 => X"0E4800A5900052C80053DD6F9415430001008AF904E064A15488843130702E30",
            INIT_RAM_06 => X"632A011E72100B51258B1386A01942B3E2752A88B1512113ADD884A728022520",
            INIT_RAM_07 => X"94D0610C90D3139308577F7DF7DFFD7D77D7D7D7B09D662C44E042016A34A5A5",
            INIT_RAM_08 => X"100A20E2329899264DB12640914A9A1A0AD12849213C34483941842470D94715",
            INIT_RAM_09 => X"73A672C32A6DB6B222ADC5ADA4C9B4090617169160842196D0135294A4408830",
            INIT_RAM_0A => X"9A664D29BB4915ADED6B79681120822548B2A92881884105B946931338C52980",
            INIT_RAM_0B => X"B18B36D8498D812B11820C6A884085A94B5909A452290C848CCC463062190881",
            INIT_RAM_0C => X"33096D1296B1336D9AD63A75DB43219210DB602CE0B6C26DB4C8582C26710D8D",
            INIT_RAM_0D => X"080993164080243534C1AC1367490201C6E1221E3B69A244DA25AC627242A356",
            INIT_RAM_0E => X"470C09763BD0641A63A211A332134D137A35E38B58270B44934A184CA0C6630E",
            INIT_RAM_0F => X"5A64EEB1B4B498063C773304E190CE3B8201D004D014D8108D80DB1C45B18221",
            INIT_RAM_10 => X"6432D72653464965A821A322B326D41CD329348948B51288122923A4A0D450DB",
            INIT_RAM_11 => X"62F4C0624E325D0249292058C6820C60220820A5DB57B56B406482A509F6308E",
            INIT_RAM_12 => X"900036CD984C2D0C0001B06C38F00C4F120832636826B5A821186176C301A180",
            INIT_RAM_13 => X"636860C5CD0C18A609265240B01A4A4846035821E2F0D4549A87A398BC30A816",
            INIT_RAM_14 => X"CE1C80100530904591803102033C7E1A9328CC025A28A47209092E580D00013A",
            INIT_RAM_15 => X"162C8E0241DC16400601DB552DA66AA5A06D0831C5E2B2C664C4989D71E87129",
            INIT_RAM_16 => X"4A16273016B0900020E265AD6B6C818483AF8C0387AEA68C711E3B013704C987",
            INIT_RAM_17 => X"C908B0204A6A1054C78B464A23249260630BAAA9B46A880268B44008656A5826",
            INIT_RAM_18 => X"827A20045690624042D4144C12A552510421954818E381128126AAC0CEE08910",
            INIT_RAM_19 => X"6D36D1AA114E1630C2CF008019224DA114E2C503163880884224C062474422B4",
            INIT_RAM_1A => X"8C6A4150942C822484091243341A2D09CAA9B8AA10A109A138AB1C570A040CC3",
            INIT_RAM_1B => X"088648764D4150052A2921CAA8A436C60269DC486BBE68B8E3486048824A6A10",
            INIT_RAM_1C => X"9364C4E56190928B59355AD369B95465995195B5B59609993356B6B0452A8505",
            INIT_RAM_1D => X"C043B70CEC889A110DE41C8072D23968105B00A407225012806D8340A6118D80",
            INIT_RAM_1E => X"122124221152906419001537129B2AD18C6142250C82424B25989619092830E1",
            INIT_RAM_1F => X"4D8910D6481B36DB6DB2D80041280201482198B6066D60430B09144009122122",
            INIT_RAM_20 => X"2D3008636DB6DB65B6D1B6D09A10D18DB4D34C0B2435851240CC13484B34B326",
            INIT_RAM_21 => X"D191B1A0606C00004D9861B6DA498024005009A680CE90A9421097620188D100",
            INIT_RAM_22 => X"DD61A4248684129D15D3A9A6F22213E6C86DB5ADA436DAD661924A02500B09A4",
            INIT_RAM_23 => X"A1B69011104104AD9C21058D9C4DB45B7B452630183603611B46D955DF2C04FF",
            INIT_RAM_24 => X"C16A089266401A340049B6C75B601B3ADAC1550268893484CCB373367293684C",
            INIT_RAM_25 => X"71D9B686C43108474EA6E5AD4C820884782380010604A000806310006219C01F",
            INIT_RAM_26 => X"2B81450A14684C0154000DAB6CD46C5B14C86889064980921864D490D8909B6C",
            INIT_RAM_27 => X"292C4E3D999A3A39C63871CE6F8E14D8D94B89248A2F9E700E0E511545045144",
            INIT_RAM_28 => X"94124C054C4CB2CE5921B0CE47F06338393876E666E7639F9D71894DA18D5087",
            INIT_RAM_29 => X"4F01C058CACA788A8A78CC9880C8135B0B24070C7231361D050ED778A2D26864",
            INIT_RAM_2A => X"65908194CD17BAF7343096678A1BF1BC1DCF78A37398DB48B6D16D36C16909A6",
            INIT_RAM_2B => X"0D340509000250898889424E9B84C899336B264D79260191089E211E93E10844",
            INIT_RAM_2C => X"9B12A444DB352C3444DB34B46C18D83086869A6014300010EC6C20DB69F62967",
            INIT_RAM_2D => X"1B62B5C6DDB1DB4360884B6C421B54523E5252936268EC37610A2265324C34C8",
            INIT_RAM_2E => X"6C4C2E1B5ED89C5A6C4F2F086CDBD1B11278DA68631B536D86031B6CEE0D8B97",
            INIT_RAM_2F => X"09B1A18D0862636C0D34988D2EDA66BB2B62676C68E8EF4DA6CD92B5764AD892",
            INIT_RAM_30 => X"6DB6DB6DB6C6276E61C31C926925424694A088209D4B6C5136D1C39045148649",
            INIT_RAM_31 => X"4AE1211075C49057122B8430233C00D20952C922419172E9243188E5C0CD8D9B",
            INIT_RAM_32 => X"9890D916891689292045165207169385BB5B4919267732AB20539C867E112227",
            INIT_RAM_33 => X"DF0C14B84B5AC312481874CA5E12D7262925A05AD9384F8D2265DB2878534690",
            INIT_RAM_34 => X"40000000049A4C31C75DEBBD3346C42C86195A0958A52109B2FB1A6804200026",
            INIT_RAM_35 => X"6118E5A0304D834BA524E6D0D8E9A60BD057921E86BC3030638EC4D0229B5000",
            INIT_RAM_36 => X"203184D6B6D87070810200C22C0040C6D042A8226892A49890ECCE4444726733",
            INIT_RAM_37 => X"700208B5810800400004400000E1C0C6630920408000C1040000880B8E00D853",
            INIT_RAM_38 => X"842011B2201903504403206A0B58C6181040202D6018C6B4210080400104A038",
            INIT_RAM_39 => X"8912616218216561165224226041805998459434EC4D261A4C9A0160724913C9",
            INIT_RAM_3A => X"9112D2D0D0D0D0CA08892C21022249040882828282828281220CE40CE11A0310",
            INIT_RAM_3B => X"C4D89CB627231A92486600ED208630B68320892C122CCA742A09A69A69480000",
            INIT_RAM_3C => X"A2C4995016B06C3C580992314B4A810B6DA2C42DB68B30D36D869B4CED9D3614",
            INIT_RAM_3D => X"2488AC825904B2083285650A4C90F14D490B8B458C30ED9364DB078A6A48585A",
            INIT_RAM_3E => X"300292984E492192312210203808438E010871C660441244464496412C82608C",
            INIT_RAM_3F => X"C000031B4EE4CA69B4514D0544810981090C989A0B596B58C040220400800818"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C639DFE78DCDA956B5AB0A2A844D4609E61664DD0124BB1DA4A52270EE1FE010",
            INIT_RAM_01 => X"14044404C6C0800D0082B1208064EE38AC49B5B20A4097FF0041859325144518",
            INIT_RAM_02 => X"8B15EF696A932C4350A25B46610C431288813999319993333B83888148D73E2D",
            INIT_RAM_03 => X"24C1082ADA40A48844349A06328B6DA0D24890D761A4DA4D369B6D949000A161",
            INIT_RAM_04 => X"1DB23F66861FB64C1000454150B43F0000B55605FDDFD2430000000040001011",
            INIT_RAM_05 => X"17E04103FC2081FE10810082101041C0200000180A40202010008812508E0211",
            INIT_RAM_06 => X"00841080D0421C3A12002048040AC0083508840402C2048010302103F024081C",
            INIT_RAM_07 => X"3BC5A6D5EFA96EC936820280A8A28A802802A802D20820009210084387402A12",
            INIT_RAM_08 => X"C9183253683101505AE24C816BB123232122421FB3942142E11F435BD257BD31",
            INIT_RAM_09 => X"C0A9C214C3EFBCFD4512A9CE0A6324FD9787EBD1C48ECD6B38650C610811029C",
            INIT_RAM_0A => X"D7D39BBD52B4C9CE7CE49F1466C419E0A6B157410728951A6CA9DC7A919E9391",
            INIT_RAM_0B => X"E30C286E7200A1A32F6ABB9125540086318C0094F67B937B590C82D06088482E",
            INIT_RAM_0C => X"4FF51F2A72A2DC10610B810201A65614550EC7DAD0D38950C90A77D9C892D130",
            INIT_RAM_0D => X"5E3837524744D14F696A5697939792935C8AB5AFDE67E6550DD4AD45B49C9854",
            INIT_RAM_0E => X"9AE1D6D594A708D0AF0A662EB1EC766E4BE4BE895AE52955914E2A954CA5C638",
            INIT_RAM_0F => X"216EC462265123880CF403FF8221367BFFB5479947994EDA6AA6B6289E9D64F9",
            INIT_RAM_10 => X"614DAED1CAF7765E4F723BBD2F398E7F45D251379392D1177BF1FB3B3D27F932",
            INIT_RAM_11 => X"937D6893CFE15A0497FAE56D2693956A82BFF0C3A6264A462E7BCF674670B1F9",
            INIT_RAM_12 => X"B874E5D794874A3DCF129A59B12224B675924D04912C62533CD7592D840962B8",
            INIT_RAM_13 => X"B4A8F126D71C24C7125CF5CADA25FEB96B44D93D565729A8416755529549134C",
            INIT_RAM_14 => X"39CF3EE3EA5D688C82A28144F96A96A4A554568DA8D349D3DF9B1DA04B1E369E",
            INIT_RAM_15 => X"79FE31AD17217B16F0F43288F912D11FE27938F32CB6B1C8F7ABD054CB2ACCAB",
            INIT_RAM_16 => X"B46833B7E7382D9F78D8D94A52816E416CFE836EA2F5DD764CD67BE9E4FA3460",
            INIT_RAM_17 => X"0EC78CDEB844EFA31E2A323CEB23B1EFEB3D14128291343AA3D126796291B1AA",
            INIT_RAM_18 => X"C993DE1C85F989BBC88865B16D1A2DA499E58A3622802043CED111311A082604",
            INIT_RAM_19 => X"57430A449FBB30836A172FC8604E50C9FBB21CF450B9FC27E4E548939A7BE42F",
            INIT_RAM_1A => X"69019E8289D6B28FCB8197BBD1A8D04F48E62A8A38BF9609E98835451F23304F",
            INIT_RAM_1B => X"BFEBBFC91617311E8CF3F54DEB1CFB7FFC1210229010D24B821898673DB945E7",
            INIT_RAM_1C => X"67AA58FA1A1F6D318E1214B1B8EF8523322CA2E2E223E557B50B2B2F898DCB88",
            INIT_RAM_1D => X"451E48A517209DFFD67FEFC1C255E12B6D8DA34BE1674DBA6E46D5A348AFA39B",
            INIT_RAM_1E => X"E84E84D6239772B626B522C40AA411479CE752E715687DB55A4A21A1F6D8B122",
            INIT_RAM_1F => X"9754FCAB2F845B6DB6E473FDBFBDCF3D5CF28F747C36D6E736F3E7B7F1204E84",
            INIT_RAM_20 => X"1A9518D56FBADF7D9E739E799B339738E38E39345B2B791945962E6CE45E45CB",
            INIT_RAM_21 => X"266BB186C50793C90874AAD3E8F4E04C1C3093BEE1633198E6718BE50DB9AD11",
            INIT_RAM_22 => X"DD5574478EE470A93E8D145114467527C8CF39CFA4679CE7AC9669B74D94D44C",
            INIT_RAM_23 => X"E37C9132145145A9CAB5B36B02CF6F5ED49366729D3EA60A1284B5F9A02804FA",
            INIT_RAM_24 => X"BF87ED16CCC073BD88FF2CA02081230104100626CEB26696AA3B8AAEF997E8F6",
            INIT_RAM_25 => X"B2EF36CECC739CEA3451094B58E014187EC01E44110007910080401E01000F1F",
            INIT_RAM_26 => X"514156A455294C814000892A4B99EC7B08ECF6ADD6FF229231408C9199999F6C",
            INIT_RAM_27 => X"6318C210E88808104208208421081090D0420DB68823AAA40FFAEAB82FFAE804",
            INIT_RAM_28 => X"FD324CD8875AF36F55BBFEF727A2E73030306666666663199B031B1FE318318C",
            INIT_RAM_29 => X"EAB5AA8FD7D71BD5D51BCF9689AE4D7B032DCE6A62E1745B103FDF3CD9926892",
            INIT_RAM_2A => X"6771339CC1F31A63BC3D26739A07B9B5A22E514496B9F9DE73FC8E38E1D91145",
            INIT_RAM_2B => X"A9E7EC288B68B905FE18E82D322EB7B46FD30D9B8FFE169C0ADFA38EFBFB9CED",
            INIT_RAM_2C => X"BF2460F6FC69CCE0F6FC6F70CB7F96FFBCBFF7FFF7AD3323AFFCFB1FD17E4E5B",
            INIT_RAM_2D => X"BFC62CAFF9F9F24644140F5AE73F19E7DFC7C7DBE77EFCE4DF9814FBF8DCE7A2",
            INIT_RAM_2E => X"E8D8BD1FFCD5D46AEAEA35792E5CB3FFEBEE3ECCEEB7DB7DF66B5A4E7A391952",
            INIT_RAM_2F => X"19EB33599DD6476CFD75D1EFE7B7569467C6E7D8D8F8D2F9FCAD46696E59F1DF",
            INIT_RAM_30 => X"4B65B6592CACEDCAC79A18A3EA098BCFDEF2D8A942235AE7EFDD29C9EE7BF2C9",
            INIT_RAM_31 => X"63EB7BA6C7DDB55B628FA470CB3C44D23D5ADB6F64972A5B6F9F1549B5995976",
            INIT_RAM_32 => X"F5CBFF99E799E7BDB5E6D96FBDFABACCFAA609CBBD2B7FFB795E908CCA390CAC",
            INIT_RAM_33 => X"F39CF6C51B94A8BAFE4D9D12694DAED1ED8D4694B8A5385DF9327C49A53BEDD2",
            INIT_RAM_34 => X"600000000C8A4656C76CED9DD354ACBE8FFA54EA5E7394B1F9BF33CE446210C7",
            INIT_RAM_35 => X"653BD1382A0B45996C6DCFF4915F3822751FB6338CDE323246A78CD13AB255AD",
            INIT_RAM_36 => X"306313DEF5D614158B14D7DAAA3D68E7C5853386CA166D921570F766CEB87FB1",
            INIT_RAM_37 => X"23210529514B860618688B005A448CA5C638E6C58B26CD34C30D1162DCD9DD24",
            INIT_RAM_38 => X"15BD296A0B0E6D4B0161EDE97AD4A572CDC1A0CA58318CE7085B8341B4151C91",
            INIT_RAM_39 => X"891AE744B8FDE6E25E68AC582C978939F8B79AB57CBD271A4E3A6D37295564CF",
            INIT_RAM_3A => X"8DDBD1D1D1D3D1C626ED9CE159BB671C689888888888888EBBCE7DCE7E414152",
            INIT_RAM_3B => X"77BFEA6FFE8A339BC8E296D3264CE6748BE2229C6BB7CDF4701D75D75DEFC5D6",
            INIT_RAM_3C => X"F3D096D0FB294AB8F5094AE53DBEA0A6CB36729B2CD9E1BACB0DD65ACB59644D",
            INIT_RAM_3D => X"B26EECB7D96FB2DE0285250A5C97D19F59AAEDDFB8E24B42D0B23E8CBADFF06E",
            INIT_RAM_3E => X"B35B9EF94721A8D9B5C478E35EDCEB96DB9D72DE29B4D937665FF65BECB7E36D",
            INIT_RAM_3F => X"08C35E367D336514428A722996E3CFE79F97D5D4D2956F79CA651B91A2D32319"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"21094FF5E657C804844D3A04DD4A6EC942CA740152AE1A8F24205D8F01E01F9B",
            INIT_RAM_01 => X"847E580A290B51A1D719288A5BA4AEA8B4C86A22521BD2AA0A44848D1B7DE884",
            INIT_RAM_02 => X"4026B400E25AC3F913118B2426E7F90CAAD7777757777777777C9D4204114B08",
            INIT_RAM_03 => X"C12A49056C9FC9AEEB6DBCF34D74B2592C977D74BE596DB2C92D926927DACD61",
            INIT_RAM_04 => X"347BD261430964A8AB451014555510100082A000A2A22024FFFFFFFFBFFF1B42",
            INIT_RAM_05 => X"E81FBEFC03DF7E01EF7EFF7DDFDF7D3FDFFFFFE7F5BFDFBFDFFEF7EDAF71FDEF",
            INIT_RAM_06 => X"FF7BEF7E57BDE3C5EDEBDFB7FBF53FF7CAF77BFBF53DFB77EFCFDEFC0FDBF7E3",
            INIT_RAM_07 => X"50E2A10280C3068D080282AA00A80AAA8002AAA82DF75FBF6DEEF7BC78BF95ED",
            INIT_RAM_08 => X"143198C2281025996E301718050A46060E5561896115B8C06F033802DF450DF2",
            INIT_RAM_09 => X"DE82DE017A4926D5E6B46528D30DB42906179091428415105A11CA5293807030",
            INIT_RAM_0A => X"FBFB0DADDB06B5ACFD6939A3129E327C103EF5E871E32C60AB7A95531CD8E188",
            INIT_RAM_0B => X"31C871014452C90383A2DC8A545BFE61094BFE4C120984103E6A1A57685A3806",
            INIT_RAM_0C => X"07030D3E12180524AA52AE5C253398D9D623E12CE498C0E2122C5D2C93181382",
            INIT_RAM_0D => X"B51C7D93E234A6467B42241BA7010B4DCCC0747EF9E1B76E207C8530312F82C3",
            INIT_RAM_0E => X"2F22696EB9CB11CD34D08AB59EA8E0966864C6F99C75FD05D9EB04229494C259",
            INIT_RAM_0F => X"475053A2B68A440BB9A49F05BE070CD3829129022902208CA8C2EB0624450129",
            INIT_RAM_10 => X"7807DB776FD2C1642820E962B5EAD43E28248A0924DE06843227E9F0A0165053",
            INIT_RAM_11 => X"285040286CFACCC1252AA1C84488373C440920C6CB5C176B416082A60BFC1FB0",
            INIT_RAM_12 => X"E6842761FA30AC7EE88C406C38702603201517252826B4BAA152693AD181A050",
            INIT_RAM_13 => X"2118205085080A1D0486554390094AA8CA0150877E611D5D8E15CDCF9801AA34",
            INIT_RAM_14 => X"7C5C410C3082C048F28099010B2FDA0A88868400052092DF0F8FB40C0D040128",
            INIT_RAM_15 => X"040D10468E1002815C081B552DA6AAA5A06D8C717CC4F6C2ED429AB95FA05D61",
            INIT_RAM_16 => X"02038632B6B41269896C6DAD6B3896A0960EF816FB368215E11CD314660EFDCC",
            INIT_RAM_17 => X"793044110F7B18552A43D3C979F5FAE2E280EFA4642A480B140A51883D8A18B1",
            INIT_RAM_18 => X"C6D7000456F8C24D40F6161812A55A5D4220F74210BE08168177AA508F800980",
            INIT_RAM_19 => X"760890A9110AF04BDE0780820511621100AE0C0DF03C800941366028DAE4A2B7",
            INIT_RAM_1A => X"E23A605032D9C7448031228B0A05228979606F92912500512F94BFC94A0802E7",
            INIT_RAM_1B => X"C8024B805501D000E22161782197224401ABF750285365BBBA882609C2073B18",
            INIT_RAM_1C => X"3210C6C1043200594BBDD291A8C9763D336D94B4B4B25BB931D2B2B2D862C594",
            INIT_RAM_1D => X"515C050C646AF11004C09800DE416F21022100020B22525291708500034B2D08",
            INIT_RAM_1E => X"42B42C8E045250A6006915FDD6006A23084363758210C8008418B243200870A9",
            INIT_RAM_1F => X"D58281D05C59524924964A01210807086C705C240684614202842409055AB42B",
            INIT_RAM_20 => X"0C310861C9239247145114529A1A918CB2CB290080758DD61154036C6B56B56A",
            INIT_RAM_21 => X"C207B1A27C71D226B6B3B10805020814021005A6884A580C4358CA60C5874068",
            INIT_RAM_22 => X"3F8E1C1A8354309D1EF5EDF7A2A253A6C86184206430C21065B1CA4A52602B83",
            INIT_RAM_23 => X"309490C7082082D6188436A5103092E2F3489421DBB3A2411B46CA217F8007FD",
            INIT_RAM_24 => X"40780732EEC03D22042F964FDF7EDC7EFBEFF9E174EB640910C42443C6604421",
            INIT_RAM_25 => X"A2A9248484210839D3B784A55DCFEBE6013FE03BEEFFF80EFF7FBFE07EFFF000",
            INIT_RAM_26 => X"FEABEAEFBF961C0155507D836590ED1B435B28DA4624EA921D33E39030907648",
            INIT_RAM_27 => X"BDEF7BDE8EEFEFDF7BEFBEF7BDEFDEDE9F7BE924EFBF24DAF5B5EFBEBAAAEAAE",
            INIT_RAM_28 => X"A0D24C6D7D618E8EA369679D5618C21FDFDFBBBBBBBBBDEEEDFDEDE93DEFDEF7",
            INIT_RAM_29 => X"A8541781707016707016602AC65A35294365C40BC0599E1D875AA6A0A6DB4C69",
            INIT_RAM_2A => X"BCB0D0E6622080103124B085136F75FB9FED69A53B104C25984B30C11F290492",
            INIT_RAM_2B => X"071CF8E284EC5889DEEB3BCCB301D9B16629AC588B2C143A70CF1B87D9B1086A",
            INIT_RAM_2C => X"A216882395550858239554A039107221C3C44A402211001199D84120A9802524",
            INIT_RAM_2D => X"026070C083079A6243EBF8844A00C4427C80806540A0E876E8F08E4D12A85C4A",
            INIT_RAM_2E => X"3C0C0280022891C01448E0385CB9D00126E8896861004E49240A11B4CF1901A3",
            INIT_RAM_2F => X"02106083082341C81924900D2294D7916141162C22A28706A3AF1615235810F2",
            INIT_RAM_30 => X"6FB7DB6DB6DEC6EC6302700D346444C884250862BDDC844300694236CCB09649",
            INIT_RAM_31 => X"C48093A6ED05092736920C34EAB000D21D3A28AF60B336652ABB1148B09DCDFB",
            INIT_RAM_32 => X"889603329B329B0840CC32C26D7312BE8F00B898D5628550F4ABD8A6ED1AAF8E",
            INIT_RAM_33 => X"BA486928595ADD05011A325A8A37DB77D22CAC5ACE28DE86246CC16A28C44891",
            INIT_RAM_34 => X"C00000000EA3505B82794F29EA49446160FB4AEB4B084A532CD21A6939094A4C",
            INIT_RAM_35 => X"EF79CFB527194509A6B784B5F96DB497212496190530B8B8C36884D028D21B18",
            INIT_RAM_36 => X"CF318D84269A525089158D7B59E09494E2D28A2E78B2659ED369D655FDB2EB08",
            INIT_RAM_37 => X"790698B5A9091D5D34C4440048F1E484C21871CBC71D9A69A698889EF98950D3",
            INIT_RAM_38 => X"0FB42F2F0E8AD264E1D15A4C921084DB9A4361AD60108421002186C348CBEC3C",
            INIT_RAM_39 => X"306363440F2A333C2337B6377468F6CC0F08CDE748A9A4B248D352E966B11ACB",
            INIT_RAM_3A => X"F44670707070707A1A2367B5A688DB8E2AB5C5C5C5C5C5C4331EE71EEFF07B04",
            INIT_RAM_3B => X"D5EDECFB7B3718C6E83668EDB5B6B59EC030D447834666A5529DB69A6843455D",
            INIT_RAM_3C => X"A24A3A84F1766E6CB8E3A3B498A997536DB40D4DB6D034DB6DA6DB6E7DCFB630",
            INIT_RAM_3D => X"0DA206680CD019A1F6042CC9C633D714CF7EF9249C70FDC771DB1EB8A67BFAC9",
            INIT_RAM_3E => X"66342A98EEDE15B6B362336D524839E549073CAB66F386D11330033406683DE3",
            INIT_RAM_3F => X"71A6373B56EDDB7DEC59552589A30A9319149C9D8B5AC21085D2CB6759ACCEF3"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"7BDB5FEECE1FCD4E52EFB9AF0D2786E4AA5F7755F9AF8FDDB6BD000000000034",
            INIT_RAM_01 => X"D57C1D8A3983AAF5D3B9BDC77BADF63A9D9CBF2496D2FAAA2C01A5EFDF7DFDEF",
            INIT_RAM_02 => X"5AA0B6690C02EE2257BBDF6CAF8A225EEA1D5FFD5FFFFFF777C927EF6ED675A9",
            INIT_RAM_03 => X"004924A049201240600008049008001201041008040040009009248248001525",
            INIT_RAM_04 => X"4C7AED94679241E6AB14000500111F8A98882A80A20A80040000000000000208",
            INIT_RAM_05 => X"0000000000000000000000001010410000000000000000201000800000000000",
            INIT_RAM_06 => X"0000000050000000000000000000000000000000000000000000000000000000",
            INIT_RAM_07 => X"0AC5150082DAC648A802A80000AAA0000002AAAA800000000000000000000000",
            INIT_RAM_08 => X"57D2AEBCDA6D4150528A8685482500A0A91BB522427BAAB4B655BD526F90A6E7",
            INIT_RAM_09 => X"6F286CA41492494873C6AE72924A4A8254EF802AB529465245556739CADB5EA7",
            INIT_RAM_0A => X"6DBDA6D60CA02E72939C2404A8C6BA8A84A554550BAAA55432A820E5AD79D055",
            INIT_RAM_0B => X"8A5548415010AAAAA04AA325095400B39DEC00034DA654021D0F85EF5D56B64B",
            INIT_RAM_0C => X"50A472FCACAA90924738274E000742141508942295522A90800AA42202AA1450",
            INIT_RAM_0D => X"50A2A45497492542000A10A4A484D493956A1819641059B309796B552C072B95",
            INIT_RAM_0E => X"8CA80869252342D40542A048A50C641292A92B32528E72552514A120116B35AD",
            INIT_RAM_0F => X"A95095484940003DAB682CA0DDAA85B450250068006809DD729765AA80165402",
            INIT_RAM_10 => X"4A5338B700B5B490969A1AD84E512B5E08200249001295548D845A4A5A490D04",
            INIT_RAM_11 => X"A5420AA5097A92B4248495214955595D76A0071E20AE829CEA5A6A4A75E5267A",
            INIT_RAM_12 => X"25AF59152584928D105292B2A54AAA85A42443718749CE14AAE4BD59653E4E03",
            INIT_RAM_13 => X"0506874AA0D2A951D081092A42A92125285525559C964A0A554E565725D6548B",
            INIT_RAM_14 => X"B2920241001243A92C7BAEF502F3E5A16000A0AA01248064A2525109F270E921",
            INIT_RAM_15 => X"96AD5A4EAB5A52A506A944FF82549FF4CBB2528BB9348D2A932A7AA6EE4AED4B",
            INIT_RAM_16 => X"014254A419CB4800079796739C8F401A435F3D437CC150599555B452A956EDD6",
            INIT_RAM_17 => X"B504135241554A4B8F0AA4A80A4A25DADAE15550BB8503D2A0105D254AA50528",
            INIT_RAM_18 => X"296C85EBA9257D412AABA90DD250AA4970952AA1FFDF5E957537FF0FFDD7556A",
            INIT_RAM_19 => X"8242EE14252CE5439CA4AA2BA142508252CCA946E5252B5414250AA52D909D49",
            INIT_RAM_1A => X"4855492AA86C69E92A5C74A242410093B3CA373AAFD05412773C3B9D54AAD0A8",
            INIT_RAM_1B => X"BC9240D254A525D0BFDA9FB68A56F13EFC05BB5485555076DBA681AA5249554A",
            INIT_RAM_1C => X"0F009494A0A8500CE5BFE7249244294A44816A8A8AAA04442D2A4A4821513242",
            INIT_RAM_1D => X"9F7696AB540AA579249492BD6CB536CA40002A82D255A84D4250142A80084A52",
            INIT_RAM_1E => X"0AA0A900A0284A84A10BAAEED4A95500D6B4948A5012A1400016AA0A8506EDCF",
            INIT_RAM_1F => X"D59492C85C95524924954A86A0D6E9A8B69A160B5680E434A1A01B002152A0AA",
            INIT_RAM_20 => X"DDAFD6E412482490492A49256CA52A52492493A800B39D55DFD5A1B6B753756A",
            INIT_RAM_21 => X"40004E54E9502C99209BDB800004975354AF504927490552B4A52095296909D5",
            INIT_RAM_22 => X"5D249152284954AFAF3E7DF7F776D5FB12965EF6094B2F7B49253509A8090082",
            INIT_RAM_23 => X"9A016D002CB2CB24927392B14A808240E5041B5AA548F4EBA4E9211CAA8400FD",
            INIT_RAM_24 => X"000005A4FF9F7D2C2AA0596000000000000000B4748DAE502288A88AC0005680",
            INIT_RAM_25 => X"080249292B4A528CF9F7EE728DC0000000000000000000000000000000000000",
            INIT_RAM_26 => X"00410005101006FEAAAAA25494A512A4AA0824A904A4B72DBA55D82545650492",
            INIT_RAM_27 => X"2108421088880810420820842108109090420924882305101544514014150151",
            INIT_RAM_28 => X"8045B2A2A05492494922483955AA949010102222222221088901090921081084",
            INIT_RAM_29 => X"3D394A100B0B570B09574A4B2A0B40426A496B7FB292415255B8D6E1C22492A4",
            INIT_RAM_2A => X"248D5A934A0BDD7B9849DB3654EEF5FF3FEB7CF1BBA50824100824904922D6DB",
            INIT_RAM_2B => X"25960948284EA56522AAA2AB55A8DBAD58852B5616D9040F7169D6D76D9AD6B0",
            INIT_RAM_2C => X"A1A956A56D53B686A56D565EAC7B58F6DADE25EFD9CE3BAAD7B693AD85DB7394",
            INIT_RAM_2D => X"A9B5DB6A6AD56DB5B4000404B5A97FB5FB3535093524B69BB293A9E38286960A",
            INIT_RAM_2E => X"2686800000097BB684BDDB4556AD6A87B5B6E036B52921B6DB71EC00BDA6D6ED",
            INIT_RAM_2F => X"D0121A90D6A5B536A6596D4B882417255C1425A6A080A580322E55C24A5705DB",
            INIT_RAM_30 => X"34DA6924DB66D3B6B4DFECA92086E8126B5A1288000004B6C2494A003B6D64B6",
            INIT_RAM_31 => X"4A6A12F7B4F9235674A9F9777AADF524A66CA209B5245CB4482C446135269689",
            INIT_RAM_32 => X"696840ED60ED60D6853B6DB586ECAF796B612296114AC112980BEEAEB7AC2FAB",
            INIT_RAM_33 => X"2482B03554672128249528550A4338B7602A10E729291E94B054A1542908306A",
            INIT_RAM_34 => X"00000000031D8E0CB68BD17A0E904A84121AA10AA010843A4824A49212108469",
            INIT_RAM_35 => X"947390D84A525852C9492927EC36DAE1AF5324AD6EB0BABA9748292571768D29",
            INIT_RAM_36 => X"248A506B5964E6E5224010428DA50129C50944A9E6A489788C1D2155DD0A90AA",
            INIT_RAM_37 => X"4BA8A1CE52521151450EE8001295292914A608303181228A28A1DD03761D2541",
            INIT_RAM_38 => X"543B0248A0D00B52151A416A44A5295A9D144A339AA5294AAD522894255186A5",
            INIT_RAM_39 => X"5CB894D2A84524219242C9524EA482494864901A3636130D26AC61044A49691C",
            INIT_RAM_3A => X"96EA4D4D4D4D4D49AB75048842DD4051CABA2A2A2A2A2A2B2AE298E2955F024A",
            INIT_RAM_3B => X"1A66469999A0A52A16A584944611CE912A8AA32432A5483742E249249294B0A2",
            INIT_RAM_3C => X"5C90AC1FC458B4F6AD0AD29942122028B25880A2C9620A2CB251659292524950",
            INIT_RAM_3D => X"84B754A429485290BCF9B9F394A5E65192777279228A92559524AF320C93BF93",
            INIT_RAM_3E => X"58400925094129282D3744100C92AA5592554AB248F5C25BAA500A5214A421EB",
            INIT_RAM_3F => X"422840A491CF9F7DF0F3878E109A7220424121201CE435AD6A01238524920A4C"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_funcl
