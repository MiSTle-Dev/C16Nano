--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10.03 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Thu May 15 13:06:34 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM_funch is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(13 downto 0)
    );
end Gowin_pROM_funch;

architecture Behavioral of Gowin_pROM_funch is

    signal prom_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    dout(0) <= prom_inst_0_DO_o(0);
    prom_inst_0_dout_w(30 downto 0) <= prom_inst_0_DO_o(31 downto 1) ;
    dout(1) <= prom_inst_1_DO_o(0);
    prom_inst_1_dout_w(30 downto 0) <= prom_inst_1_DO_o(31 downto 1) ;
    dout(2) <= prom_inst_2_DO_o(0);
    prom_inst_2_dout_w(30 downto 0) <= prom_inst_2_DO_o(31 downto 1) ;
    dout(3) <= prom_inst_3_DO_o(0);
    prom_inst_3_dout_w(30 downto 0) <= prom_inst_3_DO_o(31 downto 1) ;
    dout(4) <= prom_inst_4_DO_o(0);
    prom_inst_4_dout_w(30 downto 0) <= prom_inst_4_DO_o(31 downto 1) ;
    dout(5) <= prom_inst_5_DO_o(0);
    prom_inst_5_dout_w(30 downto 0) <= prom_inst_5_DO_o(31 downto 1) ;
    dout(6) <= prom_inst_6_DO_o(0);
    prom_inst_6_dout_w(30 downto 0) <= prom_inst_6_DO_o(31 downto 1) ;
    dout(7) <= prom_inst_7_DO_o(0);
    prom_inst_7_dout_w(30 downto 0) <= prom_inst_7_DO_o(31 downto 1) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"4F580638656FAF3DB1A468C13B1BAB57FBDABF6A55A5552EB078601E4C0AA7AC",
            INIT_RAM_01 => X"AF017C272F7EDF52B5A700D46F9BFBE8AA5CE0914F76FEDFC25F69C020933195",
            INIT_RAM_02 => X"0836334557272051295A59EF91A539D7DF9F29C8C4A542BFC393AEBBCB4408BC",
            INIT_RAM_03 => X"97B7FE265F39E6A125EB6F9280B4994AF55EF7491187BE72D62D03E010DD7E95",
            INIT_RAM_04 => X"F46BFEDFDB8A41E15EC99F3AF498E1AE074E43FBAFF7EBA24479EDE78B3AF26C",
            INIT_RAM_05 => X"04E262238B9052083681A04E447023BAE4082347B80E8A0983391A078A7BBFD7",
            INIT_RAM_06 => X"89796A884A03EC708C561B1580511BEB974AD7AC9DD65768073DEEFF2FF7D469",
            INIT_RAM_07 => X"812C46CB0C034C6AD3418B0500C062436100D2C5500D028A63FBDCFDC87A193F",
            INIT_RAM_08 => X"6936ABFD9750556CC3DB8BCB5D77C2F801B0A6225546650D802896534A6399A6",
            INIT_RAM_09 => X"4197B891456A341943F27DC4CA2C5ACBA861486907616CCABEF36F5A4A7EE6FD",
            INIT_RAM_0A => X"103DEB9FD51D0FFD7A23B6DD4EBF1623F6DD4ED5161013FAAABAAEEAFA425FC3",
            INIT_RAM_0B => X"2F1DBF615EB983EA9E27404B10C414C89937739AFC8ADFA8B077216A9FA0B63E",
            INIT_RAM_0C => X"8DBAF5AB56AD59B316C533B595F25AD22192192DA81D8247AC7648B813B5D878",
            INIT_RAM_0D => X"99DAA8F45AD22192192FA012F590096BCCFA2753D10CED574790096218218288",
            INIT_RAM_0E => X"197BED84D053096C6A15E4D127C914C753141A48867A19AA6804BE150AF00B62",
            INIT_RAM_0F => X"57E885BFB697D611F93B91F84EE1246A7AFB4BB93F82D0345568ACD2A42542D1",
            INIT_RAM_10 => X"62F7E5B090FBFDA44E0D7DFDF8FDF8FB5DD39DB19DB0849B635E5575C41189D3",
            INIT_RAM_11 => X"1893760084490A406506E18E148BF06F64487F6248E388EFFEDDF887C5F087C5",
            INIT_RAM_12 => X"694034A01A502D29B1A5005A500D280694C27A5BBBF0722458AA1690B20B9090",
            INIT_RAM_13 => X"8EBF4000348000F48000F481AA4120E4FED38001A49686AB1D2D0D563835A282",
            INIT_RAM_14 => X"12F771F63027C4A9CC9480033084071145F813E254E6D29001912115CFA620E7",
            INIT_RAM_15 => X"6E8020A50BB501AA40000416945FF76A1D7474E7D583E591EB07A96E04512EE0",
            INIT_RAM_16 => X"D4CB27F056943BF5FCBF5FCFC1B97B7A523FAB4A76FB685FEAE8F16849240128",
            INIT_RAM_17 => X"4634821E90D21643A0104B6A63AD75FA50162626F4D4A56DF463EC5FC06837BE",
            INIT_RAM_18 => X"F35C996A2DDFA1FFBA58F4640A460CF88D7CF3D99B67D15081A04C0C7E18F80B",
            INIT_RAM_19 => X"0201A47952D29390FBFA60FDF97982E0F1A49A0B17348B1CB9A998BE66FA1F51",
            INIT_RAM_1A => X"63806F5134EC1CD1824510E404694232A11CF18AF576B916084979ADD6EF2108",
            INIT_RAM_1B => X"8A389011484A15E9F2A3884CD1B89E6231C094D02C62C096009696A28926AD6E",
            INIT_RAM_1C => X"98B41515F6FC04B2240A10B2A4CEA654AB2684566AA00A65AB68D93795EC95D4",
            INIT_RAM_1D => X"4A24D404540489981268B88114D601970CA344D579598865B6A002DA4ADD6FC2",
            INIT_RAM_1E => X"E3B159A290BCC9317E5D90884089A30A8580E0DC1B810E4EC87E296A3C5F69D1",
            INIT_RAM_1F => X"002A914D282C8F193EAAA34C1A494597A96C8C8597F377950352A66563B577D5",
            INIT_RAM_20 => X"AF3D6BD91BD97DC8A95C9EDD8B14FB52088724CD8A5D640B13449620480A6C07",
            INIT_RAM_21 => X"DBDA30D8FBB4BEEA9E2EB4FACDAB5CDBB7A7CF950A1C5544D510E921B04161E6",
            INIT_RAM_22 => X"29AF03B500287B5D7EA7AA42441D0E9F1DE5950902DA0AC1E826AAB75BDBEBF4",
            INIT_RAM_23 => X"B8D11F92BE62930A5744E48D5DAA5D0AAB82430CB0C0241042481F0032B8A507",
            INIT_RAM_24 => X"055300EE200E30320D16B4E2205A655B4353AD40DC2C864F1AA50E45363EB0C5",
            INIT_RAM_25 => X"82BA7AC0E66189310AAE1ADCDCCB3B93179333EFD2AF8BCA4F08B1590A3189B7",
            INIT_RAM_26 => X"D413317AECA9E1A7EB90590512EA39E2B4982A5875810D57B3632685A4E9AAB6",
            INIT_RAM_27 => X"FBAE6F12A2592320918C84BB65B5A20E8AFDBDEB3E5EF59F652F5DAE5D5AC2BD",
            INIT_RAM_28 => X"A42915D782A3C56E5D3D8AF6250096DA4B15F96566BE2AEC04D71B993B3CBF70",
            INIT_RAM_29 => X"EBD2D02D16425A0161A0BD02F491642C20FB727445A4015569300D2495425157",
            INIT_RAM_2A => X"8B649523832A8034A9A0192FDBFD9ED3FBC9F93B3675FEDF2FA7FE93F23E4D95",
            INIT_RAM_2B => X"84D8BA4F9E0595EBFEDAFD2DFE1908A234AEA2F5D2EC2C9E209250BB751353CC",
            INIT_RAM_2C => X"F53DD3F7748680F8BD5BFBDDCBF54AF6CE49B729649E5F662E6E4DFDA36AEE09",
            INIT_RAM_2D => X"6A69009A1653E4064A3B4B68148594F920053891701826E65D0D76594BACF1D4",
            INIT_RAM_2E => X"954A0ED28DD0B952AD36CFFDA33BFB7047B3EFD4D6520F79AD93A3122140C947",
            INIT_RAM_2F => X"B3F5FA5EBBAF47B06FB46D7DBC48923EEAD8D9F2C4FAEBEF549D797AE8349058",
            INIT_RAM_30 => X"DA496B4A46918D2A17314FE0808B04845469E1DA4F7B2A0000D00149145874A5",
            INIT_RAM_31 => X"F40B888296B698C0C0C16EC050F85C76465B5CB36EDC28A8EF547F0949CD6295",
            INIT_RAM_32 => X"DF5326C0B36039AF68EF3ECC7256B1EEE7F6DAF27476D7B6FE9722B9598160C2",
            INIT_RAM_33 => X"1EFD427E27E4812D22F7ED822260EE714D611D72A3E2764E6BC56F87A3F23B46",
            INIT_RAM_34 => X"B4F1BCDA358690A4575F86BC5A0FB46F2FF74DB3D72205194C0B62D108B4E78E",
            INIT_RAM_35 => X"64D80C9429136630C69A50D09D8065A02A1C118D3662C6C69A81F81A3E49CF6E",
            INIT_RAM_36 => X"5A1E5B50AB1F4340A3B81C3729450D82BAFD0804C4A01399209A2EF7AF2DD02A",
            INIT_RAM_37 => X"A49B89825620F879740B902E4947F5DB6735DFE88748D81A08748D86C25B12DA",
            INIT_RAM_38 => X"A215432499124D821D126C36287A59756CC94F570EAD16528885DAC8D24F2593",
            INIT_RAM_39 => X"DDC39AFFF77ACAA355AC8460125043F7CB10C5CF1673E08EF436676276633201",
            INIT_RAM_3A => X"E3DBF8A16BEE25ADCD21A190C4890D0C1011DA6CB41363274085A1AA94B4811E",
            INIT_RAM_3B => X"000000004E30019EDF6FF3D90D5EA82BDAF600161792365CD4EB08C93DA8516F",
            INIT_RAM_3C => X"00000000FFFFFF7F00000000FFFFFFFD00000000FFFFFF7F00000000FFFFFFFD",
            INIT_RAM_3D => X"00000000FFFFFFFF00000000FFFFFFFD00000000FFFFFF7F00000000FFFFFFFD",
            INIT_RAM_3E => X"00000000FFFFFFFF00000000FFFFFFFD00000000FFFFFF7F00000000FFFFFFFD",
            INIT_RAM_3F => X"60000000FFFFFF7F00000000FFFFFFFD00000000FFFFFFFF00000000FFFFFFFF"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0410422824260C051D5B43405334008050A4021680400202D048240424800208",
            INIT_RAM_01 => X"0D98A080000D44042108280800040D12040824A526D8452074A02A8144804900",
            INIT_RAM_02 => X"4804009022010F24021004AA5D004009005088A0C1009184A044102081B71620",
            INIT_RAM_03 => X"86194B24A0908C9002019004082100048A915204050924D51003846000A32002",
            INIT_RAM_04 => X"09A4C308A420244210480910A408A0059216A021865A9152482200B0810C4240",
            INIT_RAM_05 => X"4C400104A8AE2228052802240402111040411444000008908016001909B4C209",
            INIT_RAM_06 => X"2D142E4620122AD8640025A15B09D61148040016C209420B4C92004300210480",
            INIT_RAM_07 => X"001048042C042C00030214200500905495009100B01012DB489148908A445905",
            INIT_RAM_08 => X"80D0804BA417403714856D182043644004445010012884A22024A84081452209",
            INIT_RAM_09 => X"A9C6A4EB512D2A9C0B0101271A8140A033322604401754D20092E928A8482A19",
            INIT_RAM_0A => X"3605100C612806C18190CA82004C81930A8200EA80A4A4200004004300B4A012",
            INIT_RAM_0B => X"840814090A10B5026A0083043120000A1420A01DDA48184800A36D0918401614",
            INIT_RAM_0C => X"56F4A88D1B264502650C4A12901188AC624E24C240C0DB2841000E14DA12A52E",
            INIT_RAM_0D => X"2509410C88AC6A4EA4C000D908016CD10D409A40231284A02091608625E25A85",
            INIT_RAM_0E => X"4F400BB006806CD5408582048048312AD4A055C1A906245000B6428842C03286",
            INIT_RAM_0F => X"CB4A0C9B3E159610412010614C08BD424850D55905284091D30A071200008840",
            INIT_RAM_10 => X"2806509262CD44C5A20D0910B258A0D2108B516C59F8109A634A400009A40217",
            INIT_RAM_11 => X"1C4537506C3D827870AA65C506D411020530652C330D330CA26800019DB8061D",
            INIT_RAM_12 => X"493D249E924F69270924D6924F2927A4938912511100D2011011045028289CD8",
            INIT_RAM_13 => X"0B522534A534D2A534D2250804882C64150869A529042011CA0040239635005B",
            INIT_RAM_14 => X"48A2182002249424842D9802022005404A01024A024295B30143082481095045",
            INIT_RAM_15 => X"E4252904C08108068B4D252493008280202A284A848890248911040210000421",
            INIT_RAM_16 => X"341320A58848106405012C4802100C20DB485249A91FC8610004800821260400",
            INIT_RAM_17 => X"212920A9B43FD5D03F09201B09658836A8B2F0E0080F08D0421286A042409052",
            INIT_RAM_18 => X"261236949362130B1B426362104610DD0C550B44C16D02004B361A42A5868480",
            INIT_RAM_19 => X"141421184981945853430B520D0D111510962923016A3441635F42688126B464",
            INIT_RAM_1A => X"C13D204DE13624092207B19775312128034A0BE100D3429AA440A04128904850",
            INIT_RAM_1B => X"32914B02845A36C108291525AAA5AD150490A2041B548804040401084D29262A",
            INIT_RAM_1C => X"9420040D126110208106302081002462CE8C208AC0068892110D02C820486044",
            INIT_RAM_1D => X"5AEB352D352CA4B0B2C46A0B621214D29B065A60843427DA6C1338A55A112192",
            INIT_RAM_1E => X"B55A14410914352493484516C58DAD508912508701510816FA93284216084206",
            INIT_RAM_1F => X"530008282228A806A8D36348527BA684C49B5B120168834D06F1A6188C40A0A0",
            INIT_RAM_20 => X"84240A4A2D0225209342306941E540B68254A0C92C1165024300842519488118",
            INIT_RAM_21 => X"7EF233ECA138E847141D2FD4AAC389E5C6AFCF7F5F218A092628A001240845A8",
            INIT_RAM_22 => X"00003020CD050083001084D32D08A1306110512230015AA94A639A7F4E9D4BB9",
            INIT_RAM_23 => X"A067143450C89E650D91AFA604A142640694D24D24DB6924D8D2132500214961",
            INIT_RAM_24 => X"509420A88408814290140202905090528201018C20241150A13E446D9C08A0A6",
            INIT_RAM_25 => X"56A15650818026140B401F8CDE9A159FB1DFAEA6FFA4703C92A0222960291260",
            INIT_RAM_26 => X"2D468495120D289110B48B48201431B8B6EA0488D8DAD69208B1B1108530B000",
            INIT_RAM_27 => X"02010588F904885A4422514E904009B4A58C522096AD184312B01AA112D4B929",
            INIT_RAM_28 => X"0310B22039FA92D186936C4D5F7245B5B0D894D89369AC016280A18440000004",
            INIT_RAM_29 => X"16240740452F40AC04416405880052F00A0040981C0849862C8206209B220801",
            INIT_RAM_2A => X"50011354586C01123006A0218C209B424989A1644810C30936849A1262C88202",
            INIT_RAM_2B => X"4F84368C416C96080808080B3690041241A81020A0DA6509081484A620BE0606",
            INIT_RAM_2C => X"D8C208B6590B10B0A18D325B7A44DF4C6B6C3EC016C0180102092830D802D94C",
            INIT_RAM_2D => X"DC40405861A6064090B6F14202C86981B3098C080B05882410CF5B9634D244F7",
            INIT_RAM_2E => X"98812DA7581845326582908098106186B404042054D8690CA02A0B20B2081216",
            INIT_RAM_2F => X"09000502853626CB6212251284121120800548C0A45404200D86B58AD0190065",
            INIT_RAM_30 => X"B0E2C14010145842181918321A903D3422C305B75820B12D28614B04BA009A13",
            INIT_RAM_31 => X"02020539D104434B4B44D25A00018051968083104103642D0436901324283039",
            INIT_RAM_32 => X"088081B20619861241868209080DA61044DA00B5A50C625369001088152B1B28",
            INIT_RAM_33 => X"C400322C26405A01AC1A105292D3029A052D654C20C2600106960C6A152C8630",
            INIT_RAM_34 => X"4906622590A80C02C804B104C960030806120923465890B4B9260DAE43426DB6",
            INIT_RAM_35 => X"A92313634008CC451DF0424943448042364994988CC5011DF182020C90531010",
            INIT_RAM_36 => X"108088323158DA0D8051C20A054009624310D369911646400D201340C4B129C5",
            INIT_RAM_37 => X"C6400FB468AD0D8583C40E107AC89004008341804581A11004581A44093649B1",
            INIT_RAM_38 => X"46964B10900848011624D22001020210C05BE85862181800D434300863605610",
            INIT_RAM_39 => X"00984180A2042B519836854C106026D620804108A2426D280024004015901606",
            INIT_RAM_3A => X"58611610900001000D515118C0428A891445A587CB100541482896C082925091",
            INIT_RAM_3B => X"000000360541B2420CB09145612C641020226D60C28DC4C30B18449A0016D106",
            INIT_RAM_3C => X"00000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3D => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3E => X"00000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3F => X"70000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_2: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"C3484C10473DAA6CA92A4A00333A03C1E9DEAF7E45AD7500E170458C68A661A4",
            INIT_RAM_01 => X"8D71CDE3637FDBF18C63781C0FBADB6A8A71AF817FB7DAF7FCFF61CE19F40D4C",
            INIT_RAM_02 => X"0C0207545C2D60531AD6D16319E35B16F6CD6500FC65413DA3F196AFCF551F8D",
            INIT_RAM_03 => X"35F6DD1EDDADEABB072F79F189AC1B19462887C5348410775C1D8DC0581E5F95",
            INIT_RAM_04 => X"BD6DF6DBDE8150810E619728E0B040EB150867DEFDB7A8A42D51FF570E1EF125",
            INIT_RAM_05 => X"4994EED4A28402645E7C1608395CEA98A2C05096F80C08808BB61EDB0B7DB6D7",
            INIT_RAM_06 => X"4A181566013F226245B4092C127D9B69972ADFE49516536BEB2DA0BF0A52F483",
            INIT_RAM_07 => X"1111C8440C340C0A1B1A54056D00A1458C62911970D03ED048E9D4EF9FB08A63",
            INIT_RAM_08 => X"E9F6E3DB251671ED937AEB6FAD5F5220B55081017058A16A000AA8475C11A209",
            INIT_RAM_09 => X"B5C7ABA4516AEB5D6BF6715D22A95E4E29592B256D522F939EBFCB7AEF7A2EFD",
            INIT_RAM_0A => X"8092ABBEF508DFBD5A59A8450E5A825AA8450EAA83C182FA0AAA0AE3B074DD0E",
            INIT_RAM_0B => X"3B94FDE112218FE0FC0F030F84C002CF9F114395F84A55481423802A55400712",
            INIT_RAM_0C => X"DE394466CC891871F3E0329465E3C27F019899E7EB9F193EF87F54E8CA94D554",
            INIT_RAM_0D => X"194A65F8C27F019899E7AEC9DFD764EAE7F83F47F80CA5370F0061F0998198CD",
            INIT_RAM_0E => X"765A7B74779664EC2C15F5C18FC380CF13354F8C067819F80BB2763E0AF9F9F0",
            INIT_RAM_0F => X"EB20A7DF3FA3971049209048C82F99035A31DB6A63421430967AA2E205AD0E4A",
            INIT_RAM_10 => X"FA97FC3BE0DFCFE1B72E5D39F0F9E0C2D5CB956C1DFC18F6F29E94558165415F",
            INIT_RAM_11 => X"14D5AD08A45D067053AB516A8E9BB9AF21B17F7C330C330DE7FCA2A3096AA449",
            INIT_RAM_12 => X"5056282B1415AA0B5141635415AA0AE505AB34179798BD24103B84082073BCD0",
            INIT_RAM_13 => X"87BEC49AA81A6AA81A6A2800D81006398C4234D540440366D48006CDA929B5CC",
            INIT_RAM_14 => X"6E5749722103000B0C1489012B029161EDD081800586A29188E0B5BD628631A2",
            INIT_RAM_15 => X"5E216501402180DE11A6ACA5055BC728947170E721CDCC16039B930638092E82",
            INIT_RAM_16 => X"76D14C68421219F564895EAE61B77FF8DA77B282DEF6D07FFDA6C02401F3110A",
            INIT_RAM_17 => X"2D0E288FE4BFA7D23B09690B6A65C47CF4B2767649CE9CFCBE50F5DD30489232",
            INIT_RAM_18 => X"6D02ADEAF7D6A29C961B904F38013C042C1D589FF92BC6F1C2A116CA3F96E487",
            INIT_RAM_19 => X"104415175F4317DCF89A6FFFF54982E1B982B06A80542A74FBBFD2F0EFC57D57",
            INIT_RAM_1A => X"B23D7973C1FAAAC621420177C9F9615E015B9F6BFFBEFF182E594AB452290D51",
            INIT_RAM_1B => X"B9A9DA09751C3FE07A1A99EF220D2E741734B186DD410C080008C78E0C8AEF06",
            INIT_RAM_1C => X"6047031877FC44403040204071C83672E5EB45CEA9B010F69B49CADE31657CC6",
            INIT_RAM_1D => X"56DFE80BE80BBF282EB9D3C2F01DD765D685FFFCE7AFADB6DE9128AD739DEFD0",
            INIT_RAM_1E => X"1B2D1020EAEA5B696D94A432100B4A0A5A16B54B4AD09637F2AD308D2C1720C7",
            INIT_RAM_1F => X"D25E38709ECB279FCBF782FE5FFFD2F7E5B6D696F2FFF3F955A3AE35AAD553BB",
            INIT_RAM_20 => X"3E3F03FE9D8FF1AAE670FBEFEBD57FE088EBE2F6042072045B960827D348A855",
            INIT_RAM_21 => X"90FBFF9FD315B4755CBD57F55C21F8C99EF882828A7DF567C2994CB2C16885CE",
            INIT_RAM_22 => X"782F7AF59C7C7BFC5EE5AA073594A87970D8ACB60BE80A24C9538A3F378FC617",
            INIT_RAM_23 => X"382522B1E8EA5C0F4F55FDBF07B9708E2F01804284280508884A54ED1AFB8221",
            INIT_RAM_24 => X"94276068C128C85514239E84A08EB448D500E485D778165CB86D0C10AF343952",
            INIT_RAM_25 => X"C28330D6A3F1CF1685E7199FA88CE95BFF35FA37D5DAF27E7C240339E60A06D4",
            INIT_RAM_26 => X"F9C5E7E9FF8A75C76872CF2DD62631B83FFC2A7474821515F3E5219C619178FA",
            INIT_RAM_27 => X"52ABEB8A5FDFAE7BF50F85F5FC55AFBABF7E7FFBF73BF5F3DC2E173E1FA87395",
            INIT_RAM_28 => X"A231B8B5B35157FFDFFECE7A7E72D3FFFB9CF5FCFFDF4EA54A948B1568540A14",
            INIT_RAM_29 => X"B718B48B55FF593F0D407081EA495FF813941288552960822B0602C4885C41B4",
            INIT_RAM_2A => X"807D1BC41BA4603611E0A05E73CF8B416508B51D286F3CF3328651132A562A14",
            INIT_RAM_2B => X"0FC9BACE0061917BFA7B9C6B784A4192088B8279F0FC0CB04592202FCC3F3F15",
            INIT_RAM_2C => X"FCFFFF57BED7817EBDCFFB9FF3F6FFFE53583FA32487DE820B0A597DE01AFE29",
            INIT_RAM_2D => X"FEE1E0B133E71452323FF2EF15C2F9C528AD6A0010082A31944E5F973FFFF7E7",
            INIT_RAM_2E => X"08880FE71CF8A1BB7F979DBDA012FBF08597FD30E4E92B41C8038A08B09A4747",
            INIT_RAM_2F => X"82F7FE7E3F58207D6EF4EC77BE745828A6047AA847E5EF6B581FF9F8F809122C",
            INIT_RAM_30 => X"FBE0E79110444D40C9144F22DAD935B0E2EF81FF5C5F11FFB8207F1FEBD034FD",
            INIT_RAM_31 => X"72829933C79352EAEAE5E73AF8F1400150C3FE995BDC25182BD42F09053BA0F9",
            INIT_RAM_32 => X"FF40A1C28701EDB405EFB6895A5E95B6A7FEDA31D5FBF397FEF10080402E728E",
            INIT_RAM_33 => X"34BDC20020079D4D4F9FFC90F0B28AAB4E057E5E2002001B6F57EF8B81F8BFF0",
            INIT_RAM_34 => X"2CB1F01B35868886E257D7FE1E2FFC092FB404A3975F9CAFB73D0B6DC2D3CB2C",
            INIT_RAM_35 => X"E9E3D7F04000EF208FF8FAD1DF80404A1811F19C8EF6968FF982FA0627DBD3FE",
            INIT_RAM_36 => X"17B233663F1FBB4D20B1C5160B555272DFFFC361D526579C0DB85FF3FF3DFDEB",
            INIT_RAM_37 => X"44820F407F8DC3C9C54A1428700FB41405B7DBEAA88DF9202A88DF884BFD7B7B",
            INIT_RAM_38 => X"A427082C2616130AA226FC427D79D877EDD3C89CAEFE1C129035FE4322484786",
            INIT_RAM_39 => X"15CADBE9C75A0990CC9FE07A812857E70A704DEA727A9D0A0026000111400447",
            INIT_RAM_3A => X"EAFBFAA5E96800000B222294A0A111140251FFE5B490C450602DE7E10411A5CB",
            INIT_RAM_3B => X"000000184940489EFF7DF22A35CB2A31AD48035294AB4216D2C4484034A0396F",
            INIT_RAM_3C => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3D => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3E => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3F => X"B0000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF"
        )
        port map (
            DO => prom_inst_2_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_3: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"31E10040456DFB1451D4750012288743B36BF5AC17F9EF24E370416248B098F0",
            INIT_RAM_01 => X"73C1F5054D4A77421185527D3EAB5FF83F064285EDBFFE738A00008D14232561",
            INIT_RAM_02 => X"A89899C1F1920C502118194440042AF5DAC24249D093EAAFE802AAFDEBD74015",
            INIT_RAM_03 => X"05B6D31C00A94A3C274BFEC362108A739B73350C4009E795501505C0204A3A4F",
            INIT_RAM_04 => X"957DBFFF4A0A19200084542B380101109500014AEDB4A20F2150A5051A2F7108",
            INIT_RAM_05 => X"806702BB2B804168892D0A4204700BA0F1493240095682A543C91CA48F6DFFF2",
            INIT_RAM_06 => X"AA2140204C644E3A08161B30B6C0013A1C2F16CC9F7C740F4A3FEC740EF5D568",
            INIT_RAM_07 => X"C02E568BE08B602248059B0014C87A5B7310E2E1C22D0AC0093A1C1D0C8A484D",
            INIT_RAM_08 => X"E81CE2FE9741717F11CE0F79D5F8F08A08B0227250577145FF8B364142621DB7",
            INIT_RAM_09 => X"FD45BFFE71EFFFD442D957FFF38C7B2AF8500A014050054BA1F7AB4B2F7AC395",
            INIT_RAM_0A => X"368B54A3706E91F7EBE2F49AF2AF81E3D49AF2F580DC907A8BA88AEBC202009F",
            INIT_RAM_0B => X"281566E26CD8290A0B00C801A465644E1C26BC9EE4CADEAB21BBED0ADEAB27D8",
            INIT_RAM_0C => X"53A3BBBB76EDD142806818A5E1181A0340C48C084A148304405050A618A58002",
            INIT_RAM_0D => X"0C528D061A0340C48C092C1888160C400A4202401A06294060D100348C48C285",
            INIT_RAM_0E => X"3B1EF2C001570C4404A4C710008FA4628180006D03140C423B06220A52614034",
            INIT_RAM_0F => X"B4D8BB64C9A46105B05B0492924BAC2112D8C1884DA29724C672EDE4B52F7690",
            INIT_RAM_10 => X"4AA3ED3D997FBFC85F063EF9DEEFDC6D8DD1CED9CEDD8F25B39E94557759694C",
            INIT_RAM_11 => X"8D82DB81E07D8F3A3705B8CE1EC010EF48C83E734CF3CCF7DFFDA8B84C48B90C",
            INIT_RAM_12 => X"1077083B841DC20E4041D3441DA20EC107310406A6A2A408782AFE87F230EDDA",
            INIT_RAM_13 => X"0BDCA898081A60C81A604810484802B13652B4C0404601269484024D2BD9814F",
            INIT_RAM_14 => X"B7AFB4FBA5EA48E240042D1DB19A2632C002F5247120208532B970096F810008",
            INIT_RAM_15 => X"3EC92581C911104C498684B1075BD76BB5FE7FE761F7C0CBC3EFD030AF6DBF4B",
            INIT_RAM_16 => X"241909B45296337D58234E2A82245F7E9B14B883D28D927BE9A81743C8E061FA",
            INIT_RAM_17 => X"5EB7DB3EC2ED274B3895FA230EE9D13C81243020145A25B57569EF00E1012098",
            INIT_RAM_18 => X"0D4EFFA2FED2C2B4AC0294024B41CA242021C885E22B512A52E115AE7F58EA49",
            INIT_RAM_19 => X"8370FC2C7B5AC55040E30A572DD10051103123119272B97152D6DAD7B35F2DDF",
            INIT_RAM_1A => X"E5B96A5B75E82C1F8241A1F5A9ED401A835FA5ED6AF787B62E19D3E9F47A760D",
            INIT_RAM_1B => X"3BF57F081F543FADCEBF517DE3BF3B1C25FCA1D57E224A120513012AED0BED42",
            INIT_RAM_1C => X"8899354097F000980188309881523474EABB6710F332C8F7A041D3FE85C4F914",
            INIT_RAM_1D => X"56DFE82BE82BAD2CAEA0528AD45F8725DFB7F6D9EFEDAFFEFF3228ED73DDE9C4",
            INIT_RAM_1E => X"799C7C823E78FFF9FFDDF5CC160B4F60A49EFE5FD391664FF0FF11323C1CC305",
            INIT_RAM_1F => X"A434E80522EF88AE1CB682FE1FFF45E7EFBE9EDEB6DFC6FDC7E43C56AB586666",
            INIT_RAM_20 => X"BFAD6ADA8BDFFDFCAF56FFDB4AD4DFF080F3E4E4F84D7C0983819227BB48B456",
            INIT_RAM_21 => X"10D335998032E0DBF0568EDA2B01A0891E0AA88022B755675082610C9011254A",
            INIT_RAM_22 => X"11827B79101412215AD5AA1F1DA12AFA742D30590BB900E16157861A020D0211",
            INIT_RAM_23 => X"BCD849032ABF942BDBFF6F3D0DAA55AAAF13C84604680518CA4A1DED2B73A622",
            INIT_RAM_24 => X"156743C47044715395602AACB180B5490442482D1A3CD6552AFF40782F0ABE45",
            INIT_RAM_25 => X"0039584CE7F7EE330AEF19D99979833111150A2EA2AAD242750B704068F18EF9",
            INIT_RAM_26 => X"F9C5F5F35FBA90F1FA424C2454DA5ADE9B652A663D830F43B813228D88E8EAEE",
            INIT_RAM_27 => X"FBEFFC1AAFF7BF7BFD0BC57AFD17FE3D2946C68EFB63477DBD8C460D4633A2AB",
            INIT_RAM_28 => X"AC4EB97BA2AAB6F5F7FF8EFF7E7ADDFDFE1DFDFDFFFE4EEFA6DF1E1DFB3C9F70",
            INIT_RAM_29 => X"EF48FC8FD3FFD03F7DF4F903FED13FF983B624B470F96B5D4BA0B50C3450DAFB",
            INIT_RAM_2A => X"D25917A282CA9876A94829D8C6DB2E85D742784D3E0C6DB66B0D758790D26F9D",
            INIT_RAM_2B => X"EFDD3C4E8A00B0FECABA376FFCD26DB6190FB4D752FF05074DB4663F1DBF6F8D",
            INIT_RAM_2C => X"B5F7DF45B6D6C56C39DFFF9FF3FDFFFEDD58BFAA748D9ECF2E47796DAA78FF69",
            INIT_RAM_2D => X"FECDC0B031E77050123FFACE15C079DC2CC37A91381C0EE79D0A76DF7FFFFFA5",
            INIT_RAM_2E => X"359B0FF7DDA9A97AF31185A5AA32DB6047000754263A4FDC493BA202307A0347",
            INIT_RAM_2F => X"B9D3193019E919B642962814A470C03AEC8CF1F013AF296A50052D40A2D730DC",
            INIT_RAM_30 => X"F9E1E4994250C460345C0460D089098022E7A1FF5D3BABFFBCD87E47F7987D9C",
            INIT_RAM_31 => X"F5E3BD8080974AC2CAC5E9282A255523424A22B15A51449887645DCA64B46279",
            INIT_RAM_32 => X"AFD5FB53DDA9FDF40DFFBEE17B7E05F7A7FEFF53E96B77B7FEE6231999AE7A8F",
            INIT_RAM_33 => X"3CB590D209A71400CF3FD5D0F2F3CEE92264727E8D209A7F7F158B0FB3F8F592",
            INIT_RAM_34 => X"D34ED46D102AB17AA56E600407418C4D3FF46083877E1D3FFC3F6FFF03F78E38",
            INIT_RAM_35 => X"45FFDFF46211AA5D7B6A78007285B4C0E827D4159AA1717B6B03F0EA4F5B9FFE",
            INIT_RAM_36 => X"1D246A542C56610481B94D37AB7D1ED3A7DE01017E02FD0444AB37F6F739EDCB",
            INIT_RAM_37 => X"A4D10A775E01D3DD571EDC7B3340FD5F47BFDFF8BF41FC7A0BB41FDA8F6D5F6A",
            INIT_RAM_38 => X"B2E599293F149E82ED26FED41015B456FB53CE96C29C16949D15BC93D24E3525",
            INIT_RAM_39 => X"9F62FB7B5DFEEAE3552FE07B2258D7E74BCE91CFF473B9AE54B2252323412295",
            INIT_RAM_3A => X"BBFFEEE77BFB31849E1293DFE6B8949C16C1FFEFF7C6B667498477AD26B7A176",
            INIT_RAM_3B => X"000000281251FA8EBEFBE4D375DEA3CA529E2677DD1FC69FF7B416D15DEAA17F",
            INIT_RAM_3C => X"00000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3D => X"00000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3E => X"00000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3F => X"A0000000FFFFFF7F00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF"
        )
        port map (
            DO => prom_inst_3_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_4: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"1921800006369D965354D58088301D0E912994A004992C01C0E0073E20180C90",
            INIT_RAM_01 => X"1F8D0040018C652509480633180C6DA508800C01A69A694A4000240A08D998B0",
            INIT_RAM_02 => X"65898928404040C210849730C242403943013148290918E6D824037139B6C100",
            INIT_RAM_03 => X"34924330226718E20419A02431290004A8954C81A28AAA020C0A000068252824",
            INIT_RAM_04 => X"5134D34D2909C1A0306C3124000001100C2601092490811B64CC8434082D6246",
            INIT_RAM_05 => X"6C0832454451134C30D0C01A00C12301D8019808018E0F08CE3F139F8D34D34A",
            INIT_RAM_06 => X"40810031081011190A0981A8000820303948D206D410416938368453486146A0",
            INIT_RAM_07 => X"18946B2538C519912E62E539814CA1C5A1878947331430136C303B1492028945",
            INIT_RAM_08 => X"3219866D8619C33649080DB006E3E002C2510888C7CAA71290384A3900882ACA",
            INIT_RAM_09 => X"698E74DB639D3498A749C3A69B14E938724648C9124492C201CA4D8D19CC0319",
            INIT_RAM_0A => X"3449100C463906930D8484822009098604822081082C2568192418C2090022D3",
            INIT_RAM_0B => X"7092C1995EB8A1010B10842022461009932088109C8C703098E6698C70309C32",
            INIT_RAM_0C => X"2054A8CD9B36611308099210CB180F00448448004C38CB0546E161C65A10A001",
            INIT_RAM_0D => X"C90803060F00448448013458A85A2C50284042680264840010D18404484C8382",
            INIT_RAM_0E => X"734C6996301B2C5286E71406108C22429901E0611214C8401D96294B73890404",
            INIT_RAM_0F => X"5385C5BFB6D9CE18F1B918F16E4D8D874810810945427834D268C0DA8E760E5D",
            INIT_RAM_10 => X"B20EDCF3F0FB5DB3FE3C9B77BBDDA8E2718777223FB23CDA633A30C6230B8193",
            INIT_RAM_11 => X"91896449824082464112C518804449E633F8EDEE3BCF3BCFAED883C3CDB3C74D",
            INIT_RAM_12 => X"654432A259512CA981952259512CA88654C0195A1A09983268627A63D2049109",
            INIT_RAM_13 => X"8B5B0090721241B212413211B050A12514012483900C46C338108D8676339089",
            INIT_RAM_14 => X"7E0E82699C3B4619444424656F88CCF2222E1DA30CA2C884C6F0409313110020",
            INIT_RAM_15 => X"6C048535004311B6510490A65449862552E1E2C65F8FC467BF1FC11B9C249D38",
            INIT_RAM_16 => X"325128A8010951450155A948225B4920C118D32A6312664924840731C99189E8",
            INIT_RAM_17 => X"0024454890240C40E4012080284128A404208292A18958905002922293000542",
            INIT_RAM_18 => X"B41F2496924A52121922432DB89C3AB015872E24084907C986363001A4028006",
            INIT_RAM_19 => X"8D3368DB4906CD724A1928542D05695B48412C1300C964C94652464E9D3CA4CC",
            INIT_RAM_1A => X"9C23A0C50324E284112497149323B34C104B013582D206D4E0C986C361309236",
            INIT_RAM_1B => X"6496489ABC8126C2884927A65054CD920E50C408F109404B9CCA8C0C08983439",
            INIT_RAM_1C => X"AA541D925A48625122A40651A39076418ADC06C2911411D21929864C366D405C",
            INIT_RAM_1D => X"830903C102C0B67702D3677061200E0E520C5B4884B4E492490131B646313519",
            INIT_RAM_1E => X"0542325979306C07B618CF3A8B0418B39E81C94C876F153C81B664AAF23AC48E",
            INIT_RAM_1F => X"B49421D4E8001A695A8A40487249358C86DB3B3B636D22600C8D025ACD690000",
            INIT_RAM_20 => X"7736176DAFCDBBE3D063DF7DB9366D040D8B11968B2AC5E5721C4A46800DD2BA",
            INIT_RAM_21 => X"35C6D0AAB4592D4011C670D9CAD502A54757F57DFD60888985AD58E2D1C4A33C",
            INIT_RAM_22 => X"C058696822C2C002420C66826028F120C01C863F2286739852065F66AE2316BA",
            INIT_RAM_23 => X"E751AF2430CC536D8D19A4E42461C26C2664120D20DA682619D07300296F68E1",
            INIT_RAM_24 => X"D08E4D51E193F1C410CDAA1983369098DA092D6148413138F124812434296175",
            INIT_RAM_25 => X"9CE714D183619C8FE0C60EAEAA0E559D555962270F00525E9838D3098B569248",
            INIT_RAM_26 => X"A30C8C80121D6DA13126D26DA0066B61649A26DB189AC6129805B59833E920A1",
            INIT_RAM_27 => X"66CD310C0924D9CE4ED26A409046DD31A1091024D488126A5861B0E1B0C104C3",
            INIT_RAM_28 => X"14C6716B04043881269A4C68C8C769212498D690934D1CD6919A6D19B0DB6CDF",
            INIT_RAM_29 => X"C626DA6D8926902433B3691DB490926D821A5BB46D702D4509A0DD08D640936B",
            INIT_RAM_2A => X"DA699F083B4A19B469B669A529A6DE9AFF6DF9ADB4529A69AF37B7DBF35B4D1A",
            INIT_RAM_2B => X"6D8D36CD30E9B069A86911CDB6DA69A6899DA44133DA4D024DA426760D362684",
            INIT_RAM_2C => X"90924904D33A2FA6F38DB73B676FDB6C686D368036D69B43324369249211DB6D",
            INIT_RAM_2D => X"DB6DB39831B624381976DA6D8CC06D8933118C041B0DB1A4D808D27424D26C8C",
            INIT_RAM_2E => X"14D23DB698C083F3ED1684849252493631911434CCC349059D0733033067032E",
            INIT_RAM_2F => X"114630E1F1AD05BA4A51A3D0846098208492449BA2842118CD0423078375A359",
            INIT_RAM_30 => X"B0C4CB320C93206F143860209199098032C31FB61829A924625648A496661810",
            INIT_RAM_31 => X"62060D04899653474744D609858184CD82C803114842650D252694D245283037",
            INIT_RAM_32 => X"0985CB8356A1B4D009B49B65E8EC14D3069B6DA58D08631B4D000944B719E708",
            INIT_RAM_33 => X"C484235A35A413209C1210D1D1D343C32CE9ECCC35A35A6D364C38620D22C612",
            INIT_RAM_34 => X"51424124D6185359852DA4449B4B584134D864132E6C1876D8361DB607630C30",
            INIT_RAM_35 => X"11BB7B63040488D3492051006306A06C2C059610C8894949200F6C3A0E5B3F6C",
            INIT_RAM_36 => X"3001041860B008241093041258E3B6C3021049259882660085A0924084E32799",
            INIT_RAM_37 => X"A4D2C810CC3D858D068C1B304480905A469B6D338B45B62838B45B6A0DB66DB0",
            INIT_RAM_38 => X"880C41266F13378E2D36DB5042C20110C04768314A59711AC2143067D2625CCF",
            INIT_RAM_39 => X"991269B1046C4E491064864CC8D446CE18860118B046293814600120CD80080C",
            INIT_RAM_3A => X"CB4D32D9B1B013102CCACAF8C1865654080BB6C6D112518DC00DB68046529F97",
            INIT_RAM_3B => X"000000206AD1B61349249AB8290848294B5049C33A69205A6A0A320A58C459B4",
            INIT_RAM_3C => X"00000000FFFFFFFF80000000FFFFFFFF00000000FFFFFFFF80000000FFFFFFFF",
            INIT_RAM_3D => X"00000000FFFFFF7F80000000FFFFFFFF00000000FFFFFFFF80000000FFFFFFFF",
            INIT_RAM_3E => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF80000000FFFFFFFF",
            INIT_RAM_3F => X"F0000000FFFFFF7F00000000FFFFFFFE00000000FFFFFFFF80000000FFFFFFFF"
        )
        port map (
            DO => prom_inst_4_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_5: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"41CA1186BC6CEA0821204836E4F4D9ECE3CEE7399EFFBFB48C46BD0E9740A0F5",
            INIT_RAM_01 => X"236716FD89EB557BDFF5815CAECE79222A6595EB3CF3CF7B8133B371E6998201",
            INIT_RAM_02 => X"96525311592CF6DFFDFFEB5379FFEC5D53B3290A2ED32D35A7FAD3A9CD4D3FD6",
            INIT_RAM_03 => X"6EBAEDC3BB694BA3EC4D62BA69FEAC48130265FB3A528B6400C0300F8300AB4C",
            INIT_RAM_04 => X"D7AEB2CB39C340AE88D635E793461A22FDBB894AA79EF26196D38C4C68CA5489",
            INIT_RAM_05 => X"9320CA06447CB59728AB83CA92DDAE34B07A88266F4CBE157A357293B9E7965A",
            INIT_RAM_06 => X"B0987E4089C2596E4328537EB6B39A2335B9328DAC54C69B5A658955B8C558DE",
            INIT_RAM_07 => X"B05D8D9727A6C60E11D3377747D9CF46ECCE85DD4E9B572590E337D5204D7DCD",
            INIT_RAM_08 => X"3C94B35A4C6359AD671899412750DCCDBA76220A5F4EDD13A0686E8D7629F36D",
            INIT_RAM_09 => X"27252A81C94AA877367A65554EE2CF4CAEF3DE7FC3FE9A2622AA994A5A589297",
            INIT_RAM_0A => X"49B022C25D0D619D0E98A114CB0AEE8A2914EBAAEE96DD4CCE74CF8E2CC9332A",
            INIT_RAM_0B => X"7273F3E9BBBAD18E4DC13982C99D0D7B76C512F5857891607836937891687419",
            INIT_RAM_0C => X"50001354CD53321C28B26739032C14159B29B20A70192DEDCEE480CB6F39BD17",
            INIT_RAM_0D => X"339C892B14159B21B289C36FB921B7D8946313B0AC99CE446166305932132EE5",
            INIT_RAM_0E => X"F5FCEF9FA820B7DA837B481CC174C993264682B66C99B263B0DBED49BDA69459",
            INIT_RAM_0F => X"C72DA4BBFF91DE71773371744CD45753EC9F777DCDB0D11D7DEFC8F36CA66DE1",
            INIT_RAM_10 => X"6E26F9A753F25FE33E4C1763389D29DAD393916D59F97C92653D36DC54136B37",
            INIT_RAM_11 => X"F7616D378AD270D7D8C2D36B61376FA663AA6F48E269A27F2FF98E95576E94D7",
            INIT_RAM_12 => X"E6D9736CF9B67CDB8F9B5CB9B65CDB3E6DC7F9BA3A24B2622B2E68D342C51724",
            INIT_RAM_13 => X"529753E773679CB3679C337F6DAEDDE73611CF399B253DB39E427B673CF3CEB2",
            INIT_RAM_14 => X"6FB5BE4FF78D5739577FF6CE4FAD88F73BBBC6AB9CABCFFE9772CE5563DCC610",
            INIT_RAM_15 => X"EC927E4B6D09FF69AE79DFCE6DEF1C765B55C7ACDD6D5AB6FABAF6AED8FEEB7E",
            INIT_RAM_16 => X"C9A7B9B6118DB3531337399894BACB2924D6A736CE76E7CB28899E698B1D28EA",
            INIT_RAM_17 => X"77D8F64B3F6D8CBD27FFF614DDB319ABBA49CD8DBF1B339157BD88BBDEDE4DCD",
            INIT_RAM_18 => X"F473E49B924E26323B8E45F966B4A1B57F9D3EA514B91CA772AA97762DFD8FFC",
            INIT_RAM_19 => X"2488021AC9136D9A7624BB77B71F29CB6C9BE9BF5A4C66CE56325258AB2CE55C",
            INIT_RAM_1A => X"A67B62D1CBBB2B1065CADD5F41B9C5CDD7CF2BE580D30499A9AF128944A24192",
            INIT_RAM_1B => X"38C87E2D3F292ECACC8C89BF651F0EBCEF59D070DBE5512B1C2A603CDECA3644",
            INIT_RAM_1C => X"2552EAE433C5E35518315B551BF309E5F0FE8A2D926BA6F326D3976CCC36E1AF",
            INIT_RAM_1D => X"238D80F181F0F737C3C8773C644067CF7B2F5B61CEF72FDA492FF5BEE7BFA971",
            INIT_RAM_1E => X"51A8D8227E34EC85BF39D32730501E8612A3E33C33BC31ADA73F82A13BB9B467",
            INIT_RAM_1F => X"4E489733C510513ECDA2146C9BFF1FFFCEFBBB9BEF6D8676ADAED39CFCE7A6E6",
            INIT_RAM_20 => X"77F6537ECF9FBDBFE9E4FBEFDF4A7DDB78A9299287ADC37566302A9F2DB6CAD9",
            INIT_RAM_21 => X"12C210888010204010040090080100810602020A2022AA8598CB378A5702A94F",
            INIT_RAM_22 => X"0D51DCC68A8A8C45E7273973AE61A2A26739D535401CE7B27D82020242110A10",
            INIT_RAM_23 => X"7F73235A73997DB919D56FB7A5E34538F53A6CB4CB45B6D3652D9D36CE5E94BB",
            INIT_RAM_24 => X"314FDB1BE71BE35A31CA4E39A72991ED2868D21B66AE96D9F2B6F0A7FE47B31F",
            INIT_RAM_25 => X"39ED9B21F7FDEE4F45CE08888808011111110226D2F7A582596054B47245AA49",
            INIT_RAM_26 => X"79E6E6F35B288209A20920928889AF6065A0F90871272C6AAC2B6A7BA3BAA207",
            INIT_RAM_27 => X"70FDF6DDADFEFE73775B897ED94EEAE67394CF9F8A67CFC531560BD70B52F32D",
            INIT_RAM_28 => X"EA196A10F3F2D6BD5CB2B8CA4A52572F2B719C9192CA8BCEC9390E7FF21C4E02",
            INIT_RAM_29 => X"CC41FC1FF1FD6C7E55DA527179671FD64721B3DDC6A979B670DD87B398CB2510",
            INIT_RAM_2A => X"65A27AE48D1CE71B7AA17AA318E39AB379D92B277194AAAB2766FAB2566ABC79",
            INIT_RAM_2B => X"9B166B3882365AA88CAC3B9B2B2592DB56DACCE5CE95B264B6D95965B66C4568",
            INIT_RAM_2C => X"91C71C5C718AA8AB691B2AD2D257B648CFCAECCC5DAA3435E3B5A7AEA5A695BA",
            INIT_RAM_2D => X"B517A1A5594C598AA565A51D0D2A5316644D19F6ACD6613A711856167EBF5FA5",
            INIT_RAM_2E => X"592CE94D315F89EF50F866E6E5AF5D594AE88E4B031DBD1E02D6ECAECAA155AC",
            INIT_RAM_2F => X"255A52241235ACE1B39C3819C9F16EF3C96A50A44ECA39FE76E529108E1C5E66",
            INIT_RAM_30 => X"2E94B816A1B82F9E9BB6AE4F2D27E2FB8FBA3D2DB1AAF3FFB1707FD7FBA15579",
            INIT_RAM_31 => X"E477E6D16E7AEE72727E8895101B1A197D3C4627ACE4BECAD54D55249EE6EBAF",
            INIT_RAM_32 => X"091EAD6E74F777DFF735DABEEE6B6EFBFCB2EE5B339CC632CA04A205806F72DC",
            INIT_RAM_33 => X"0BCE4E6AE4E8E9FF1E32196DADAEB5B4D033707CE6AE4EADF5A4489E256F8C6F",
            INIT_RAM_34 => X"E59B643F3D5FA865E8C2188961B18EB7F5D7BBFEA4D9F125B3E4496CF2C679E7",
            INIT_RAM_35 => X"DB2AB2C4F7D8FE71EFF384BE52FCD69BB1757F790FE1C1EFF2927B8EEFEE77FC",
            INIT_RAM_36 => X"B24511B322119EFBFD9DECB368C2DAE67A31FEFF337D55FA7A725E44A5697949",
            INIT_RAM_37 => X"E96D9B2AD9D71D971C78B0E2D03AD1F8BEFACF3E8DDF2D36E89DF2C9F965CB2C",
            INIT_RAM_38 => X"ADCDBEE475723BBA274B964F880C2794E4D3D737329F96E7B9EC30C674D5A58E",
            INIT_RAM_39 => X"B3AF5D6397589375FB3EC86C84F45CA44F29AF8F1DE3C6FF7B5DB6FA896DA5E6",
            INIT_RAM_3A => X"B7CB2DE32322BA528B9697B59684B4BD7DFB2D8C96693909FEF21E8C7B7C9D1A",
            INIT_RAM_3B => X"00000015CCF5FEBAEBAEB35CC7189C339CEFB4E7B98FDFFBE7399DFCD9CBCF2C",
            INIT_RAM_3C => X"00000000FFFFFFFF00000000FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE",
            INIT_RAM_3D => X"00000000FFFFFFFF00000000FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE",
            INIT_RAM_3E => X"00000000FFFFFFFF00000000FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE",
            INIT_RAM_3F => X"F0000000FFFFFFFF00000000FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE"
        )
        port map (
            DO => prom_inst_5_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_6: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"3140E34C6E76ADB6DBDEF762D2744723932A94A48CAB3491FAFC6DE86DB098A0",
            INIT_RAM_01 => X"2DBD08A2052D6190A42A2C5229094DB21D236E97B6DA68426E22C6CF1D3BB761",
            INIT_RAM_02 => X"CD151590E89B20C10A424396DB2110506A71AF81F453B3AEF2D53AB12BB796A8",
            INIT_RAM_03 => X"169B6B7E887319AD040BA15066841025AAB54C47D3892453DE3F8FE078FF8D4E",
            INIT_RAM_04 => X"1BB6DB6D8C4178C6B40D3A758E0D31113EB4B18D66DAD15F68E6C626DDAD6247",
            INIT_RAM_05 => X"CD038F5E1545422594549E1C10C8F61593C0AA0C53381E609BE43AF21DB6DB63",
            INIT_RAM_06 => X"6EB02E7540FE1513418A0185122DB021324DD206C63B426B59A4841A48406FC6",
            INIT_RAM_07 => X"7AB97C2EE9BE08A5425F2E137D8DD976D877CB93B6F83AD34DA13386D7C2C901",
            INIT_RAM_08 => X"269992EFB63BC9778D084D02F5636805BBE208A8CF7DDDDF4FEF5C0FB083771C",
            INIT_RAM_09 => X"D9EE75FE7B9D7D9FC3D455AFB3F87A8AB5D4BA974CDA67DA02DEC90A18C8631B",
            INIT_RAM_0A => X"246B550D4CEA2695297B9C9A54E9AD7ADC9A54BFADC988485920598651A60097",
            INIT_RAM_0B => X"7DBA9127B3613807434CDD99A34CE09AB566953798D856E712AA49D856E715D6",
            INIT_RAM_0C => X"07F5A8993264CD67A668D318A2990EC74E8CE8821B9E9B7814FB5CF6DB180FAC",
            INIT_RAM_0D => X"698C048E0EC74E8CE8806EDB02D66D856E01D0F63A34C6080CDBB33468C68FC0",
            INIT_RAM_0E => X"426C4EF095D76D80F643370ECC9FA3408D0BD8ED3A04E801ABB6C073219B5334",
            INIT_RAM_0F => X"EA19AED26493253143223142C88B1DB46C16D549016057189B4FC19F05AE3862",
            INIT_RAM_10 => X"BE05D0BE489F6DFB262B3DB5E2F3B4977F8679BEF12AB2DB43BBB2CC45D1613E",
            INIT_RAM_11 => X"1ECFB78282CDB7507B9F69FC2ED11B263B215D7926186609B6F886BD89BEBE89",
            INIT_RAM_12 => X"335A99AD4CD6A66AC4CD754CD6866B5335794CCE0E19863A2166485E4076F6D8",
            INIT_RAM_13 => X"8B59ED2C59ACB1D9ACB159A4905A6A3404005962CC6F5247B8D6A48F71DA3754",
            INIT_RAM_14 => X"481700EED7FF86EF896936FE7E1DEEC1E88BFFC377C46D26F7483DAFA65B5A69",
            INIT_RAM_15 => X"3C68E98D645BA4965ACB1D3335ED8E32597365C6BDF9888C3BF36222F236EE2F",
            INIT_RAM_16 => X"B6D9202C000300698C018C4866CD6DB6DB52999ACA5FB06DB7868C2F0075E89C",
            INIT_RAM_17 => X"39AABA1DE62DAFD8FB8DB0BB6C6D8036A1867676098A18901B18C788294DB000",
            INIT_RAM_18 => X"1C3B2482924242120F36404DF035F4941CB14674FB490ED3F671B3E277C4C6C6",
            INIT_RAM_19 => X"8B62F8AD490DC269921B4B048D0C4E129AB40B41C85168D342D663CDAD342554",
            INIT_RAM_1A => X"CDBB20CBF1F6648F962D37A7E9F3B54C544B1BE582D35498661B0582C160B62D",
            INIT_RAM_1B => X"75D4EEAAB69566C30C5D25F7B0675C9E0E984533D80B0359B658AE1C2919F619",
            INIT_RAM_1C => X"E6C5A638DB68CAC4682832C4EBB100E1DEED6158D08059D3080587EC5684600E",
            INIT_RAM_1D => X"D7DFAB0BAB0B363C2CD1E382E13FCE2EDB0EBB68D63467DA69197DF7F73BB5BC",
            INIT_RAM_1E => X"2D5651C96D747D7DF7D8DAF0000B5C16FA15D70F471DF176DA77D58A769B51AE",
            INIT_RAM_1F => X"D6746DF0BBEF8E6FCA9E02EC1F7F14CEC6DB7F3F636DA26D6EECACDADD6B0080",
            INIT_RAM_20 => X"FE7613EEAD8FB1F1D763FB6DDD40EDB0DCB935F23B60F5ECDF17586FBB6EF0DE",
            INIT_RAM_21 => X"DCBBDEEEFFDFBF7FDFF7FEDFEFFDFEFDFFD7FDF57FDFF5C38CAF2CBE4375831D",
            INIT_RAM_22 => X"2414D94AA8A0A489630E700E31A8E160E31085E62BAE4B744253FBFBBBEDF3DF",
            INIT_RAM_23 => X"76C9261571DD9E2D8DBBAFBEACE1C2AC7445CB6AB6B96DACD95B3AEDA94E4AC9",
            INIT_RAM_24 => X"90AEDF1793D791CF902D2A0590B490085E2F212549543078F17E0F5C3E2BBF14",
            INIT_RAM_25 => X"92DF10D7D2CF3AAC31840EEEEFEFFDDDDDDDFBBF57FD575438EF41619BC71668",
            INIT_RAM_26 => X"3BEFCFC01B1E71E5A0E28E29D044A5286CBC703710C01430D2B1B1303B2160EB",
            INIT_RAM_27 => X"C199A18D5DC6EDFB761728E4D81CA9A135AA1C38850E1C4290389C389CA21585",
            INIT_RAM_28 => X"7E4A294A555058E1C4D3484DFEF371B9B89096D8DA695985C57059B760301820",
            INIT_RAM_29 => X"8408908933BDDA3E2F60CDB32C9B3BDDA3161F90D4AD59040F25948D9068D2CA",
            INIT_RAM_2A => X"9A5D320232C85BE4617861718DB69312490921642E98DB6D3424921242C84BB0",
            INIT_RAM_2B => X"4B09A69808C1B07D886812CB24D249260999244324B20DA24936242C892C3C87",
            INIT_RAM_2C => X"D8D34D1E9A17097463192A5652549648737C6C8426C5D2C2774259B6CA1AB24C",
            INIT_RAM_2D => X"96E9B4F2252426FC506CBBEDA7854909BCDBCE4190483DF5901EFBFE76BB56EF",
            INIT_RAM_2E => X"10926B3590BAC3264FA796968A136DA085244626ECB34D89D9066616615F8A0D",
            INIT_RAM_2F => X"106EB4793D64FC964210623294E89A71C483E7D98787B5BCE836B1E4F6512648",
            INIT_RAM_30 => X"67B19FAFCBE2A36EF3532234D192793DA69E1D65D08D21BFFAC0EFDEF3281058",
            INIT_RAM_31 => X"42F779B7CD27C767676EC7F0444D88EFA4988B125D696C7C41A606CA4C7231ED",
            INIT_RAM_32 => X"0D0CD9B74E9B269A49A6D348DCDD269A4CD34A21098C421A68C2E23318FFD74D",
            INIT_RAM_33 => X"24C617C87C87D4495C1B1891D1D343DA6EC0EEEC7C87C859A69F3E0303BCC626",
            INIT_RAM_34 => X"4B2260E57719F968E529E1141E431B42669A492625FD387EFA761FBE97636DB6",
            INIT_RAM_35 => X"B9B71F60174BDCCB0DF1B99B6B4F8249E013B738BDCF2F0DF11BE9E826D23B7C",
            INIT_RAM_36 => X"B8C044BB389CF269B4D7E69A2E58966217189349BBB4EED669307B60C673BFDF",
            INIT_RAM_37 => X"8690D9E0CD198B890D187561D11AD8D74CD369A6F90934E06F9093481DB6EDB5",
            INIT_RAM_38 => X"CEAC9A77663BB21BE4249A40A2252610D257EBB3C21A32CCC3A4307743620CEC",
            INIT_RAM_39 => X"13236DA10CC84E1B3066C0EDCAC56C851DEEDB9DE6E759BD36669248EFA48E8F",
            INIT_RAM_3A => X"D26DB48FA121A9CE79F2521792F792903EC377C59AF6AFEFE849E6853477DDF3",
            INIT_RAM_3B => X"0000002EF8C001734D34D24875AD09E1294203E2B49DD693431D36D05080BBB6",
            INIT_RAM_3C => X"00000000FFFFFFFF00000000FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE",
            INIT_RAM_3D => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3E => X"00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF",
            INIT_RAM_3F => X"B0000000FFFFFFFF00000000FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE"
        )
        port map (
            DO => prom_inst_6_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

    prom_inst_7: pROM
        generic map (
            READ_MODE => '0',
            BIT_WIDTH => 1,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"7A0A8450810903BEFBFEFF84E00E964B387039C8D1245125229086F6805ABD25",
            INIT_RAM_01 => X"827050A42A7392D294A428040212924AA275A1304924929492772758405BA0B4",
            INIT_RAM_02 => X"040202551D2D2AB5294A5A575BA56104B49AFECA25E441C923D2140A72411E90",
            INIT_RAM_03 => X"91649C02DD4AD6CD29524A12B6B5A148DF1BEB49D21DF7600000000000001791",
            INIT_RAM_04 => X"A4492492528BB96B2AA0A50CC05143BA1938C25299273AE8009729411233952E",
            INIT_RAM_05 => X"05AADCA9555554485B61FA56FABDD8B93F4AABAFE1B6AF6D0CD94765A2492494",
            INIT_RAM_06 => X"84B97FFD4F4B5D6BCBEA1B94B6F5BBCBA4024DAEC9441422D609682D0694B72B",
            INIT_RAM_07 => X"DAA7F2A9F0F950A9547CA955F45D3BF93EF7EA7A43E544410DCBA7CB016C102B",
            INIT_RAM_08 => X"4EA52492115B92494E52A240281492A8FA94AAAAB7933654FFB352AE5AAB8CB2",
            INIT_RAM_09 => X"80494828125208058492904140B09252091522A45512AA08A828A2505292A4A4",
            INIT_RAM_0A => X"4075FE1296F34920521D2ACF18520E1CAADF582A0EB49292920A9228A9D25540",
            INIT_RAM_0B => X"4A0678F64C9A82AB54150D2A13A6F5028533C6052502E577BBCC81E2E577B9E0",
            INIT_RAM_0C => X"2000DF66CD9B30802A84E8A50AA15F542F4AF4AAA4A5086AAE94252840A55D55",
            INIT_RAM_0D => X"7452AEA85F542F4AF4AA9043550821AA84AAD57AA13A29555509A54274A74BC2",
            INIT_RAM_0E => X"35129290D24821AAAA424056950013A54E95EA80BD2AF4AA2490D55521209542",
            INIT_RAM_0F => X"94BD3924C93A6954B55954B5565091A412B908302B82E72544122B3CA9C97695",
            INIT_RAM_10 => X"D9AB2DDD9B6DB27A5977ACDEDF6EDD6DEC55EEDEEEDAAF6DB4252CB110826A44",
            INIT_RAM_11 => X"444A49586AB4891514949473925BA8D97ACBB3B34CB2CCB6D9256B3AD4DB3B54",
            INIT_RAM_12 => X"2435921A890D4486BC90C2C90D4486A243432909A9A16B7A4A5992FC92A54449",
            INIT_RAM_13 => X"1CE50010521041D21041520CDE8080C0AE52A082918E7378A714E6F14A12020A",
            INIT_RAM_14 => X"B7E33AB239F2DEF6D47489795DB2EAB42DDCF96F7B6A4E91F4BA8406749D608A",
            INIT_RAM_15 => X"A2848010C9738CD8810410024336D3586C27B56B1EF6D01B7DED94072F490673",
            INIT_RAM_16 => X"4242057052952A9454AA52A281291248096721219CE4A5124A6AD17E4A97E932",
            INIT_RAM_17 => X"52949052925B0949CA94DAA1268455485C3252525456A56D2D2B2ADD490412AE",
            INIT_RAM_18 => X"5344DB686D94A9ACA8299423CAB9C82554BAD4A34926512045B02D27494A2A49",
            INIT_RAM_19 => X"0E8380A916DD0AEAA0A907A9D050EABAA9D21D2112B55AB4B5AD94B342CB5813",
            INIT_RAM_1A => X"2A8ADAB452485850942A1641524A5516943DAE5A7D2CA9A55A48572B95CAE838",
            INIT_RAM_1B => X"4A2F92A95949592A72A2BE49214952E42925705F612A5E53BF534BA68C160955",
            INIT_RAM_1C => X"4E9AAAAAA4956A99522A5299524A52152522004A2A82016CA900D4969680954E",
            INIT_RAM_1D => X"48A253A453A4094E902A94A915520B4944A904952949592596A809C914A44A5D",
            INIT_RAM_1E => X"522902ACB21EB686DB0D7ACA4894928B64A3625615BEE549235B05355A2D2549",
            INIT_RAM_1F => X"42AA95A5D50015569120A512A49243292924E4A4B496D5B4892A9267239CF777",
            INIT_RAM_20 => X"D98954929256CA4D21176592564296D04D327524F74A9BE9E8BB52A3492F3AE7",
            INIT_RAM_21 => X"108210888010204010040090080100810602022020288A24D29E75DC95B52AD2",
            INIT_RAM_22 => X"B957139DBABABB743DEB58032095DA1A95AD7FD942DC6370E822020202010210",
            INIT_RAM_23 => X"4EBB4B50CA660506D64CD9C92BDBB4069B5040200200008241012424B39CA0A3",
            INIT_RAM_24 => X"4D0B2ED775D76BB00D4A15A961286D41494A80A0B400AD65CA0940048957CE43",
            INIT_RAM_25 => X"18DC3841249072AB552908888808011111110226280008884D37B52807B5A195",
            INIT_RAM_26 => X"5ACB6B6AADBDA0825A90490482AA084D4928180B654949516143B28DFADA8AB7",
            INIT_RAM_27 => X"B566DA1656CB67BDA355AAB56D43469A1AD4A5496A52A4B52D4AA54AA54855D0",
            INIT_RAM_28 => X"BEE35B9C95550D4A8965A297B6B5A2D2D1453B6D6CB2926B554D568CDAAD56AA",
            INIT_RAM_29 => X"6B406C06DADB495B56D2B09ADA49ADB495A03F6D301C2ADB5406BBD4AD3D411C",
            INIT_RAM_2A => X"080085AAA026E9C05A3A5A8A5249A4B4925A4B4B5A252493496924B496B2A68D",
            INIT_RAM_2B => X"A6D00842AA8092A25292AD824A480002501202B4D32D04B40412424BD01B430A",
            INIT_RAM_2C => X"2565965165ACAACA4A4240E594816C96E46C896946D80404370400CB20232C2D",
            INIT_RAM_2D => X"6D04F56952D3507AA94B6807AB4AB4D4311D9C952110B5700522E4FB5B2D9329",
            INIT_RAM_2E => X"AD4832D30D016A58B4120B2B202196425202A950484802509014B52B52AF5529",
            INIT_RAM_2F => X"A0B14A954A99396824A54AA52835490A280A9529406A5AF6B0094A552AEE92B0",
            INIT_RAM_30 => X"5A6561384A13AD2FED642F50090934B0D269BE5B0D161ADBDABAB7FB6DA865ED",
            INIT_RAM_31 => X"940480950E9249E5E5E36A097574D4AAC24375A106B4048D82D64B4104A7729E",
            INIT_RAM_32 => X"F2D376C1BB60DB6D04D96CA0B6B6036DA124B452D0F794A492150C552AB795A7",
            INIT_RAM_33 => X"487BC3B2B968000497A4ED09696987690480B496BB2B96A6DB19F3A4AA4A7BD0",
            INIT_RAM_34 => X"B6D9B55B4616FB8D6E7282A80804A50519652080A9360D5B6C1B56DB05B58618",
            INIT_RAM_35 => X"D4DDADB5251D66BAE6DA4100B5A774ADDA66C60DD66AEAE6DA0D9DF6C909AC92",
            INIT_RAM_36 => X"3FB5777E4EA70804817ECB2F769AADB4A8E74924CC823308849AAC97394A5ED6",
            INIT_RAM_37 => X"6A01D2829610D0D053068C1A150F250D036D965B76D0DEDAB76D0DD6A6DB36DB",
            INIT_RAM_38 => X"6809411F594FACADDB526EB53AB8D9676D95E52504AC270ACA91DEF4B56429E9",
            INIT_RAM_39 => X"ACC1B6DAD3368DBACD592A97EAB5B32956320C521014A4B240402522AAD1284B",
            INIT_RAM_3A => X"69965A60DADA6294F3A9A9A727754D4D580A5B692C1023ABE084832840507EED",
            INIT_RAM_3B => X"0000000276B4000CB2CB35B6A452A7DAD6B525B5ADD6D04DB5A92A092D6A4859",
            INIT_RAM_3C => X"00000000FFFFFFFF00000000FFFEFFFF00000000FFFFFFFF00000000FFFEFFFF",
            INIT_RAM_3D => X"00000000FFFFFFFF00000000FFFEFFFF00000000FFFFFFFF00000000FFFEFFFE",
            INIT_RAM_3E => X"00000000FFFFFFFF00000000FFFEFFFF00000000FFFFFFFF00000000FFFEFFFF",
            INIT_RAM_3F => X"F0000000FFFFFFFF00000000FFFEFFFF00000000FFFFFFFF00000000FFFEFFFF"
        )
        port map (
            DO => prom_inst_7_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => ad(13 downto 0)
        );

end Behavioral; --Gowin_pROM_funch
