--Copyright (C)2014-2025 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.12 (64-bit)
--Part Number: GW5AT-LV60PG484AC1/I0
--Device: GW5AT-60
--Device Version: B
--Created Time: Sun Oct 19 11:39:12 2025

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_SDPB_kernal_rom_16k_gw5a is
    port (
        dout: out std_logic_vector(7 downto 0);
        clka: in std_logic;
        cea: in std_logic;
        clkb: in std_logic;
        ceb: in std_logic;
        oce: in std_logic;
        reset: in std_logic;
        ada: in std_logic_vector(13 downto 0);
        din: in std_logic_vector(7 downto 0);
        adb: in std_logic_vector(13 downto 0)
    );
end Gowin_SDPB_kernal_rom_16k_gw5a;

architecture Behavioral of Gowin_SDPB_kernal_rom_16k_gw5a is

    signal sdpb_inst_0_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_1_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_2_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_3_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_4_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_5_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_6_dout_w: std_logic_vector(30 downto 0);
    signal sdpb_inst_7_dout_w: std_logic_vector(30 downto 0);
    signal gw_gnd: std_logic;
    signal sdpb_inst_0_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_0_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_0_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_1_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_1_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_1_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_1_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_2_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_2_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_2_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_2_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_3_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_3_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_3_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_3_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_4_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_4_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_4_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_4_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_5_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_5_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_5_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_5_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_6_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_6_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_6_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_6_DO_o: std_logic_vector(31 downto 0);
    signal sdpb_inst_7_BLKSELA_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_7_BLKSELB_i: std_logic_vector(2 downto 0);
    signal sdpb_inst_7_DI_i: std_logic_vector(31 downto 0);
    signal sdpb_inst_7_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component SDPB
        generic (
            READ_MODE: in bit := '0';
            BIT_WIDTH_0: in integer :=16;
            BIT_WIDTH_1: in integer :=16;
            BLK_SEL_0: in bit_vector := "000";
            BLK_SEL_1: in bit_vector := "000";
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLKA: in std_logic;
            CEA: in std_logic;
            CLKB: in std_logic;
            CEB: in std_logic;
            OCE: in std_logic;
            RESET: in std_logic;
            BLKSELA: in std_logic_vector(2 downto 0);
            BLKSELB: in std_logic_vector(2 downto 0);
            ADA: in std_logic_vector(13 downto 0);
            DI: in std_logic_vector(31 downto 0);
            ADB: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    sdpb_inst_0_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_0_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_0_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(0);
    dout(0) <= sdpb_inst_0_DO_o(0);
    sdpb_inst_0_dout_w(30 downto 0) <= sdpb_inst_0_DO_o(31 downto 1) ;
    sdpb_inst_1_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_1_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_1_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(1);
    dout(1) <= sdpb_inst_1_DO_o(0);
    sdpb_inst_1_dout_w(30 downto 0) <= sdpb_inst_1_DO_o(31 downto 1) ;
    sdpb_inst_2_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_2_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_2_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(2);
    dout(2) <= sdpb_inst_2_DO_o(0);
    sdpb_inst_2_dout_w(30 downto 0) <= sdpb_inst_2_DO_o(31 downto 1) ;
    sdpb_inst_3_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_3_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_3_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(3);
    dout(3) <= sdpb_inst_3_DO_o(0);
    sdpb_inst_3_dout_w(30 downto 0) <= sdpb_inst_3_DO_o(31 downto 1) ;
    sdpb_inst_4_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_4_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_4_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(4);
    dout(4) <= sdpb_inst_4_DO_o(0);
    sdpb_inst_4_dout_w(30 downto 0) <= sdpb_inst_4_DO_o(31 downto 1) ;
    sdpb_inst_5_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_5_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_5_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(5);
    dout(5) <= sdpb_inst_5_DO_o(0);
    sdpb_inst_5_dout_w(30 downto 0) <= sdpb_inst_5_DO_o(31 downto 1) ;
    sdpb_inst_6_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_6_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_6_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(6);
    dout(6) <= sdpb_inst_6_DO_o(0);
    sdpb_inst_6_dout_w(30 downto 0) <= sdpb_inst_6_DO_o(31 downto 1) ;
    sdpb_inst_7_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_7_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    sdpb_inst_7_DI_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & din(7);
    dout(7) <= sdpb_inst_7_DO_o(0);
    sdpb_inst_7_dout_w(30 downto 0) <= sdpb_inst_7_DO_o(31 downto 1) ;

    sdpb_inst_0: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"D40C110B405006A5132D63084C984C4D49A9073198CC0993146331B511308188",
            INIT_RAM_01 => X"6B81059B629AD01212C243286D8A024B6C2052299EC3078504F11A2B1C10044C",
            INIT_RAM_02 => X"8D2218F22B8841860A182D003B490060DA4DB522E5D04F97414691ADA50B0E40",
            INIT_RAM_03 => X"48200D82A504444995A4A10134A1096C86248232CD40D2781E039E581330B680",
            INIT_RAM_04 => X"1844CA8C2D38B060D1C2988912E500098100101008104C0209806A25B08392B1",
            INIT_RAM_05 => X"FD6894E1DBA82A08440A21039C0300C0C0699DC7A9C476E51803542153630D80",
            INIT_RAM_06 => X"2424502290555555550B4B5D6AD50B26A24BAFB356158A0AB03418D535ED7BD2",
            INIT_RAM_07 => X"CED76D6D7BFF7AA5B4D16155555549B415BA1086FE9D7A830B8BDE27183C5B3C",
            INIT_RAM_08 => X"63ACF0A08CA20944E10A54224810AAD76B8AF016429521142A35D260A2121203",
            INIT_RAM_09 => X"819A4368BA35E9C8049D2559642425255B2BD68A4AB390B2B180B4E41668A2A0",
            INIT_RAM_0A => X"00C45245348D10402422262022262432D3962020804011A330C21023819594BB",
            INIT_RAM_0B => X"66EC549E4324BC8836A5657964F29A9A9481070422767242401201149882F014",
            INIT_RAM_0C => X"13325124226D9BD927B086282120D015088200510234A0AEE44AA0528242A106",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFF25C93F3C58AEDE480848E06B90616B5B46DD7523463144F2A",
            INIT_RAM_0E => X"FA02C3F30044C00BEF6B7BC216957D6BEED48FDD1FCC6B5A4EE3E245E413E49A",
            INIT_RAM_0F => X"FFBA034A074DF92695E0ADF7DD1EDE6AA2344D525A43243CD5C8D19E3367107A",
            INIT_RAM_10 => X"18000000000000007F0000000000000000007F00000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000100000000002000000000800000050000014000000",
            INIT_RAM_12 => X"FF0400001808000000C318000E6000FF0303C0C0001800000030060C18001818",
            INIT_RAM_13 => X"F000000F00FFE00703FF000000181818C00018F018FF01C0FFCC008001F00000",
            INIT_RAM_14 => X"18000000000000001C0000000000000000007C00000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000100000000002000000000800000050000014000000",
            INIT_RAM_16 => X"33330000180000007F0000000000000000007F00000000000000000000000018",
            INIT_RAM_17 => X"F000000F0003E00703FF000000181818C00018F018FF66C0FFCC008001F00000",
            INIT_RAM_18 => X"D1E4082A7AC26F2CDF5DA68C506400EF6B6F6FD7FAFD4404108F80FC00000002",
            INIT_RAM_19 => X"44488A448208CE9FC441C75106A21081B8268618E23D73B76DD92F91AF757EEF",
            INIT_RAM_1A => X"130402E6A48C360A48D10100A258C99091858608023AAFB72223B634032D616B",
            INIT_RAM_1B => X"2C1A94B311B8990A13690A2C88AF7D4F7D6DCA1080FCCD018300EA8A903AA3D4",
            INIT_RAM_1C => X"18F007AC64CC0BDA25A751AEEA346DA66220563342F10266B707F4E684E01420",
            INIT_RAM_1D => X"5A228B68480D365361AB8C884811ACD655DA89D4E6B4A7BFDFF767D1416280B2",
            INIT_RAM_1E => X"91096B698D84A215DA155BAE09188071D4A913D80230D0D1101EB001D8261EF4",
            INIT_RAM_1F => X"880840452D001910225AD3882B42A31A0006AC8B2C56F2B7647A2E5D220E8B40",
            INIT_RAM_20 => X"21DDF7CB9F2B751EE8DA62E1FEB4B9A388F3B370FF525CD1C479CC910F086F08",
            INIT_RAM_21 => X"FDC0E21021E01AF8612A02A843E00200026E8306004D55555A5543FDBED2E48E",
            INIT_RAM_22 => X"117B21EC80F7EDDBBF0A850487932030512443C10028041267BA1B21108440DB",
            INIT_RAM_23 => X"DFABA6F2A9218F720A37AF9C00FE057B5A57B7A1E0DB28C0E2431CC4D04877AA",
            INIT_RAM_24 => X"DD05B06A0405DD0DE01034006A07F4924124907EAED5FA8D11BFD2CE9A23BDA8",
            INIT_RAM_25 => X"833E9069C2FBF77AEDA6D3476F948629CE5369169C2FFF5D34C811048743401E",
            INIT_RAM_26 => X"C7C54154918022B02AB11840682C0350927D9EFF689F644FB5324FEF56844ABE",
            INIT_RAM_27 => X"BCE3D25A0BCA3DA127B7931013DE14E95A1AFF7ED9A5C1025F8FD12340DA5128",
            INIT_RAM_28 => X"DFAEDB472577A40282912A286818F260B0DCB3437F07A0E029AFF7EDEA95ED58",
            INIT_RAM_29 => X"12206C8499DB26F7FA8090BA80355BF7ED548A7AA50A84486A60DD97C968FEDD",
            INIT_RAM_2A => X"E40EDFBE6F7F737CBDD59F5BD1ABDB3D08A7A134690A546A0FBE4AE8411DCE01",
            INIT_RAM_2B => X"FDE7D943E244D63C6DAAAF5B4580E728B1C92AF92F6F1E647A05EA9A389A7E72",
            INIT_RAM_2C => X"B1238E95212BE25109EE25B129C146C88C42DAB5E410F0C19A1C11639A280E6E",
            INIT_RAM_2D => X"5A2164052D1010B89CB14004A0A57006DA6B505011200C8C205B0D7050C37129",
            INIT_RAM_2E => X"EF1E453FFFF8A15F8A024E465C298B5F2025C80101AD4943DEA960D0A850F7AB",
            INIT_RAM_2F => X"8522985D184008E18F2E7C7E15B44115777EFD944200FFB950FFB9516D1AAD3F",
            INIT_RAM_30 => X"2B86109680B04FBFC2025ACBE7D0A07438AD90A135A95E4222DF0D129E02B56D",
            INIT_RAM_31 => X"596FCBE4AF5C584215F4DA99EA291C24DF0A57019AE5BD5DA1988839A50CD291",
            INIT_RAM_32 => X"B54E02254B4082804AF36821120119659659C5E549C8B423E16921327C358085",
            INIT_RAM_33 => X"9697AD19972476B79FD3FB4BCAA4247023AFFC0A6925E0004390B6340296BC16",
            INIT_RAM_34 => X"32CC921E2C0E95C142B49858E89A86E4B23B5B242CA54209A6134C395508B95A",
            INIT_RAM_35 => X"04AC7942489A5088F0121A0A33B6BE9050AA7D28A257E28F01F23452E2273912",
            INIT_RAM_36 => X"F97223D4F6F949612672D052E4429937AC48AA446B13813408F528B1E3C50152",
            INIT_RAM_37 => X"FD90C063CC82D04B409184C251E04294D10240908A46A3121A4B458893C91280",
            INIT_RAM_38 => X"0000000003D7A8C1E776B7EFC025638D5111012111919191904C2257B002088C",
            INIT_RAM_39 => X"352FF340574882209A217C5018634F0C50DB921498842D4128A8B06108000000",
            INIT_RAM_3A => X"180A680806D8DC88C9ABB11928D401176D0258B982F9E73C7D7F12437C660582",
            INIT_RAM_3B => X"08241D340024C34AD28BF05807B2BF8AFF7CAFE2F899098B4E651C0899269988",
            INIT_RAM_3C => X"0925FFFFFFFE2C05850456D4A15758AAD1500A9859502BA18165305490056D40",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"61520249345249240841B24B041042617FFFFFFFFFEA29FF0000000000000000"
        )
        port map (
            DO => sdpb_inst_0_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_0_BLKSELA_i,
            BLKSELB => sdpb_inst_0_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_0_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_1: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"2C05E9B42C02449B4820EF2B260B27920524036DA4DBCA6836DB49A7864F0882",
            INIT_RAM_01 => X"842022228AA12625F55EB68892285DB49145B8C6A110693019263096C8607B93",
            INIT_RAM_02 => X"112221309AB03F5212E5C0B69210808134516944152F9454BE300809099A0553",
            INIT_RAM_03 => X"0A801210200D54088380002000003692C40C0F6D91798C91A501045064232883",
            INIT_RAM_04 => X"994000C30D12B1611081A351288804326AE5B755A8299255320A969B4A0010A8",
            INIT_RAM_05 => X"B634024356010A439056002CC499244840A8D104B015288477E3784703670182",
            INIT_RAM_06 => X"4991058410880880890096294435410A0401055221082800001471A490A62D8A",
            INIT_RAM_07 => X"9502463429ADADB0000412202202144E2410400D4990920000B8042A12801504",
            INIT_RAM_08 => X"6DAD34B3A0231CC561908404801D508A4501A4017421200754229441258FA332",
            INIT_RAM_09 => X"A50A855418316C4D08C42D496C88442C4B0816D8A025302430822606966C2D4A",
            INIT_RAM_0A => X"DC4B2EDB4C1300C06BC868DBC868D111A6886B69249B8A5533459A7D26318412",
            INIT_RAM_0B => X"2820140451A141000912981045ACA2300FE92200051100921DBF6EE0293976F3",
            INIT_RAM_0C => X"321A3A7A2D002AA850450820892E3DE24402843D4285B6C200154B840001E922",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFF4201803F5F2C96465041800521000B034548B06926120832B",
            INIT_RAM_0E => X"0399D64C38C83FE9B5B1B18307D851B6CB42AA045888429B4685269414953481",
            INIT_RAM_0F => X"FFA16A49240A452018C20026050A88029A4469BC129264133309120452A4BA54",
            INIT_RAM_10 => X"18080022004307637F1F3F0132465E063E7F7F404101007F3A01411C22367C2E",
            INIT_RAM_11 => X"0608144100003E360332397F3646403E06000800082A0000017263127F070000",
            INIT_RAM_12 => X"7F7C0000181CFF0C3CE718001F603CFF0307E0C0001800000030060C18005C18",
            INIT_RAM_13 => X"F000000F00FFE00703FF000000181818C00018F018FF03C0FFCC008001F00000",
            INIT_RAM_14 => X"1808002200447C447C1C3C202008FC1838787C00447D00787C02587F2838782E",
            INIT_RAM_15 => X"0608144100003E360332397F3646403E06000800082A0000017263127F070000",
            INIT_RAM_16 => X"99330000184307637F1F3F0132465E063E7F7F404101007F3A01411C22367C18",
            INIT_RAM_17 => X"F000000F0006E00703FF000000181818C00018F018FFCCC0FFCC008001F00000",
            INIT_RAM_18 => X"024A0032214194A28881092CBC4C940200929422901212212C1FFF0000000000",
            INIT_RAM_19 => X"240D4376582E8D28888AAB59501118575864048A0A0111A3194550C909280A41",
            INIT_RAM_1A => X"5B7030A5A89CA6420CDE75D87390CF3131B19562524044204148D42262096142",
            INIT_RAM_1B => X"20046280002A148B484298CF04063404492012940A48805285030102B2102480",
            INIT_RAM_1C => X"185822E00A014B5556215D0544B6449541075700A420147852502652C835968F",
            INIT_RAM_1D => X"7A29836900A986136051AC68608A00009504145C20C455358942030940A0E2A4",
            INIT_RAM_1E => X"23A8436C0983305868D04C36299832C4FA6C964616ED14EABE5EAEABB8CDD087",
            INIT_RAM_1F => X"348940218C221A122A10D1A812219A5900F8DB4D88BB5A61B22534101B632A6D",
            INIT_RAM_20 => X"7575F7E2F236929B622B70D57818764A9D19F86AB58C39254E8CD00154048204",
            INIT_RAM_21 => X"844280446C0B65124D41A46A582952993601B068D00666666742B36DF7D3DB3A",
            INIT_RAM_22 => X"084A11284600020400048259B0346D0582A8D833464349605406000410208840",
            INIT_RAM_23 => X"F28203431F218AA010006984BB0286AD8C60DAC1A00B01C1D6001A4400964330",
            INIT_RAM_24 => X"9A04104255850C223C00A90053442412490412420841290F9844FA859F021081",
            INIT_RAM_25 => X"A00691454A55A855452403FB4D56C65214A3691454A58AA8A4895624005BF600",
            INIT_RAM_26 => X"AC08414515E10881888000D50A80014811050869A0414020A418208446E00334",
            INIT_RAM_27 => X"8AD36397BD478955A0455604500A94D01B0369A94935794044825042E2B7504A",
            INIT_RAM_28 => X"129698452455A4000010810F5EE4AAC09C852B6B05600C4108369A943095A952",
            INIT_RAM_29 => X"C340B4A81040245142E4F6D2A884426CA6CBFE5148400002505212B136EAD56A",
            INIT_RAM_2A => X"570CFA655D2D115AD4188809408941E1AD2E23422004066A6D354A00385548ED",
            INIT_RAM_2B => X"5500280850469098B654D5880C09D68181A3B32BCC00B3374B00A29EB018376B",
            INIT_RAM_2C => X"168838244686AD844552DB1684361CC82081428064008028222015008A48230A",
            INIT_RAM_2D => X"437E98788163094A41889C43A328012112A29494C0E8E5A214221444944A96C4",
            INIT_RAM_2E => X"0000F0004808BA5405585000801428503045530A620501000005010DA2000001",
            INIT_RAM_2F => X"02005021440812858814286AB09CE200428000F57A880813400812401D1A3848",
            INIT_RAM_30 => X"42164CA68E420D3182994A800803230585000CA1516A0B0E229A2B0102241504",
            INIT_RAM_31 => X"514D50442A8884A0941116A9119C50269A2B55828A042220122B1480422A0011",
            INIT_RAM_32 => X"34167A162D0AC08B68126CB1835100480481450002000058384582342241A6C2",
            INIT_RAM_33 => X"6A5E6A490C7F6300A9766CD53420E4517A0926C82443400440C49142D7381095",
            INIT_RAM_34 => X"08936E454C65003C441C59826DDA24445B418DA9C54A20A4518187000860E011",
            INIT_RAM_35 => X"73880563509000D45870131B58297055DD2C04E84CA91047200435001412885B",
            INIT_RAM_36 => X"282114840094EA6A5504DD438903A8B41442034D4114C390110C08B26AC5281A",
            INIT_RAM_37 => X"4840BC1955A023C045D0CA6218445AD49B0256989A68A5AF13482988D00A10D8",
            INIT_RAM_38 => X"75C40001B21400187174415350041C10614151414141414150E8740522219A99",
            INIT_RAM_39 => X"8C50080B42DABA194C6815579655C456E49046A45B86C8290008B2E50231FAE4",
            INIT_RAM_3A => X"62096A76FC45544445A4189204C3E2850E484C23F0A2A0C48011AF660802BC40",
            INIT_RAM_3B => X"4D032000281398300C0510987000111118615005041D948FE302ABDCDFA7D089",
            INIT_RAM_3C => X"0101FFFFFFFF8640E0100C6040818C1461830C520CC6301A0250AE83C2100001",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"7980134DA0534D340829B24A25A2DB64FFFFFFFFFFE20DFF0000000000000000"
        )
        port map (
            DO => sdpb_inst_1_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_1_BLKSELA_i,
            BLKSELB => sdpb_inst_1_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_1_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_2: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"C84048092250C22212C4A068CD88C8CC048A25128944649200251284AB304008",
            INIT_RAM_01 => X"3114688F384C4093630C7320658132C964D44842108D128C0CD0086104010CCC",
            INIT_RAM_02 => X"8C2A18D02B984186011C6C6D81C84028502D312663F0DD8FC39621C0E5001928",
            INIT_RAM_03 => X"98C50D0528D8216A21B94200254A104003064336CD78C668DF8104482231B601",
            INIT_RAM_04 => X"8A8154504C000AF8B9A2999888220119A08100713088CD0119C2302DB313250A",
            INIT_RAM_05 => X"BF3E60488FAC1211C64C59830D0B50C04140A4B539905CF47821582658AB5428",
            INIT_RAM_06 => X"FC6CF03240473CD14503755D66635B0755699AB113048142303909C21C3D0BC1",
            INIT_RAM_07 => X"9CDF25AF2FEFEF41A085D51473CD0DBA0989B8E2F48F6853833BD6A31888171C",
            INIT_RAM_08 => X"67ACF33144220C41248A5800940888752B9A702022962282229D4AE64F3513B3",
            INIT_RAM_09 => X"AC22634C0AB12B096090E5532B0300E4535032AA4985558568C8A49C966866E7",
            INIT_RAM_0A => X"52E6DB041105921054B60225920260904B8609248208813329C390B7899DA802",
            INIT_RAM_0B => X"00A0A1019448A4D432666E0E18630C0D82C341CB001514628C3303901582C282",
            INIT_RAM_0C => X"131219341520981A302107DD821408918042481C06A96D282A8A366165904342",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFF0009282414AA938408C0442100200B53669934D3451822B23",
            INIT_RAM_0E => X"993BC2DE7B9F800F6979F9C1A7F41D6AEBF06387F44021D895A15057B5815B06",
            INIT_RAM_0F => X"FFA97A8F678ECDCA9CE7A52F0144A4D0186049D208000024DBC7CF8C62C5E849",
            INIT_RAM_10 => X"180C7F4941470F77303F7F017B6F7F0F7F7F0640633F417F7B01413E637F7E4F",
            INIT_RAM_11 => X"0F1C144100007F7F077B7D7F7F4F407F0C000800083E1C410377663A7F070000",
            INIT_RAM_12 => X"3F780000183EFF4C7E7E38003F607E03030E70C0001C00FF0030060C18007E18",
            INIT_RAM_13 => X"F000000F00C0E00703FF000000181818C00018F0180007300033008001F00000",
            INIT_RAM_14 => X"180C7F49414CFC6C303C7C64740CFC3C7C7C18406CFD007CFC035C7F6C7C7C4F",
            INIT_RAM_15 => X"0F1C144100007F7F077B7D7F7F4F407F0C000800083E1C410377663A7F070000",
            INIT_RAM_16 => X"CCCC000018470F77303F7F017B6F7F0F7F7F0640633F417F7B01413E637F7E18",
            INIT_RAM_17 => X"F000000F000CE00703FF000000181818C00018F0180099300033008001F00000",
            INIT_RAM_18 => X"D0A1503B7AE3FDEE4154A7DFFE7404B5296F39C77A278E26FC0FFFFFF8000000",
            INIT_RAM_19 => X"F50CC2E60804CB8440C38B1CA5C04C1F783E160DC1AF67D35D9139C00FE07F83",
            INIT_RAM_1A => X"13808084A488BF0BC89D67F3E3DE8F509117C7CEC2802095270BF53E2A89615B",
            INIT_RAM_1B => X"3B54B50A0A2AB54BAF7B12CF00E5ADEE156DFA100CB42A430601671483282940",
            INIT_RAM_1C => X"58B011A20A28C28203499C3AE07C6E44511385A2D439072AF743F6F7C16457F8",
            INIT_RAM_1D => X"7ACFC36C033DAE1B63EFA8EA6DC2E57208524019324845295FD72AD863C3E620",
            INIT_RAM_1E => X"81AD4BED49C6B1DDFE5C7FBE61901078FC68B79A8EA804BBBA9FEAABF8AA10AE",
            INIT_RAM_1F => X"3F4AD067CF111C151352F19A3267BA3C8002A86FAA3FDAF9F638AD149E2FE26F",
            INIT_RAM_20 => X"DB97FF0CEFD614B69439A38256EA6C62B6A511C12A7534315B5297C147423D42",
            INIT_RAM_21 => X"1586080120A02920042B92214145624892329378C627878077F74F7DDEBBA19A",
            INIT_RAM_22 => X"0252894A00522648990A110C82A10710442641502021848844CA182D72424959",
            INIT_RAM_23 => X"F4A282D38E000CC01011BF400267852BCE52BEE0C5582582A4408485544852A8",
            INIT_RAM_24 => X"9C31B36209174A4479ACACD653253BA6B26BA452CA514B0B488DB4A5B68294A0",
            INIT_RAM_25 => X"A3B2216591CE672AE490F6DACF4DA55AD2910216591C477C92082049B730A39E",
            INIT_RAM_26 => X"E52C72411DC16031E83158F0682C0294F0294A5F7C0A5005AC8805A775B322AD",
            INIT_RAM_27 => X"3EFBF98F3F77EF65FFC78A0657DCC5F2FF89D77BD490F1C005A28443E0F7144E",
            INIT_RAM_28 => X"D5A952A364440012120CA9A63CE6F142FEF1E3F3FFF7A8E3AA9D77BDF8D9CD99",
            INIT_RAM_29 => X"5251F891401306616CE6E6E4E8341BD57D555628A0811320297ADC95C85AB3D9",
            INIT_RAM_2A => X"C52AAFAC5F6E7156F59CBE5F78EF7BF9EE6F28143901455A653D28A401110A01",
            INIT_RAM_2B => X"FC3FD12BE204826DFE4ED3AF2C4AA1258849B0512D7D1C0F7384B8BEB9DC2D32",
            INIT_RAM_2C => X"A5A09298BDA58B45C014B685B04B29460A8258A82EAA10B8A22A85521187A036",
            INIT_RAM_2D => X"92D5F434A4514C52D888C446C58D6383CA28642421B14F2C6079050424B8A5A5",
            INIT_RAM_2E => X"FD16643EB2CEF015873606168A21AA96100419033CA6263C46864E5045CF11A0",
            INIT_RAM_2F => X"44B3004B142600442B2C587A9D68281505FE77C86C9F19B18F19B18918304C77",
            INIT_RAM_30 => X"01007B049CEE0F3DC1028C8B0FF1C87939AC1912101345F9169E05938C76836F",
            INIT_RAM_31 => X"534E5FADE574DEC223940132AAF608149E044229A1A01DFDE22110B3CE001A44",
            INIT_RAM_32 => X"C75DF20001280F0902D20C21000984DB6921E52048E89640C00201262F672C40",
            INIT_RAM_33 => X"99A934AE07EC52D684D2D3CE4A65AC70338FFE49000384080070A672F5B23270",
            INIT_RAM_34 => X"128A4949207AD54502B44B50E400A280BA29CFBD27054B8B6D9EFB3955F9DB67",
            INIT_RAM_35 => X"220800E00809109058020B0242AD6EBCAD5A7FE0A2D6A78400220113222D53C1",
            INIT_RAM_36 => X"5871557C322A810161224A81A04D889722AF09214293C0284891E011224417C9",
            INIT_RAM_37 => X"948282610400416040838EA058A71010594006D8004896BE5021A40A484100C5",
            INIT_RAM_38 => X"823DD55A80A8FA5E808842A8AB12E90000808C8C808080808648361180000009",
            INIT_RAM_39 => X"2C2D5A6C97020869D4082D848A26EF4E70D8A8944806A9C03C70920A09A8600B",
            INIT_RAM_3A => X"2D0F2E150444501440BA8810385C00840B559CBB57EF43687D38BE611C00C560",
            INIT_RAM_3B => X"4946796400018892248BAA4222823988B550AAA2AC1481B6DA020800B505B400",
            INIT_RAM_3C => X"B7DBFFFFFFFEEA056D0552BCB15ED4B2D0D006A8711618FB96455C73100161C0",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"B7E97497FB2C96C9F7DF6FB4FF7D2C97FFFFFFFFFFFCDBFF0000000000000000"
        )
        port map (
            DO => sdpb_inst_2_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_2_BLKSELA_i,
            BLKSELB => sdpb_inst_2_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_2_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_3: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"580CDC1B4252D0A637CB0162C91248ED1C2B11369B464092412512940BBF4228",
            INIT_RAM_01 => X"730109DB641CD213630C61636DC812C9664048298A641227EEC5CB29D1506E6E",
            INIT_RAM_02 => X"EEA05EC3C80ABDC6B0DD69DB2FAE2072EC8EB124816F1605BC95E577D501A25B",
            INIT_RAM_03 => X"48806D8605C0044B10A9890D6189196401C69BB6EF50D762DD3BEFC1BB4DC74D",
            INIT_RAM_04 => X"20109A4824415078D1219D9C0CCD311D88F90651218EEC011DC3382DB3890133",
            INIT_RAM_05 => X"ED6AF5AA41092158841AD12B10481200C829A8772C4032B057E814741181309A",
            INIT_RAM_06 => X"276FAC023612698412AC000A4C80013221B62000C4327A0C00096221776DDB50",
            INIT_RAM_07 => X"F7200D6DDB7B7A4026984C41269864014422014804010E8400AAAA0508980C30",
            INIT_RAM_08 => X"47A8F32079A705C4E0410508C820240090250942004149000980210A20000A22",
            INIT_RAM_09 => X"A9182020B820EB980C986D5B6204646D1A1176789B2271226DD024EC24E8A6C6",
            INIT_RAM_0A => X"4806DFCF3DCFE1C00093EC3D93EE60226B10E269B49B1AB22CCBB99389F908B1",
            INIT_RAM_0B => X"C46444CF074408E002876F3E50F6189F92E267E2737332344471AB8690E08045",
            INIT_RAM_0C => X"133A4C1EAA5901490280A2B8A8026044C880ECC844904D846E40927375926266",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFF56C31E4A7B162560F34FA5CDED59731F640C301E4DBA48F6A",
            INIT_RAM_0E => X"2400C6DF398D9FEAEF6B6B6035B73EEFBEDC27CFFDB9CED8DFF3C681B383C913",
            INIT_RAM_0F => X"FFAB6E87636620E6BCFFADDB40C466F820B1CF5018480030D7D0204653A60166",
            INIT_RAM_10 => X"18FE7F49414D781C1860407F49396109411C0C40367F7F084909496341490B4D",
            INIT_RAM_11 => X"59361463642449497D49451649497F45186008603E1C3E63064D0C6B14004F00",
            INIT_RAM_12 => X"1F08FF00FF7F0073663CF0007E607E03031C38C0070FE0FF0030060C18FF7F18",
            INIT_RAM_13 => X"F0001F0F00C0E00703000000FFF81FF8C0F81FF0FF000F300033008001F00000",
            INIT_RAM_14 => X"18FE7F49415CA038186040445404242444041C7F38807D04A40954444444544D",
            INIT_RAM_15 => X"59361463642449497D49451649497F45186008603E1C3E63064D0C6B14004F00",
            INIT_RAM_16 => X"66CCFF00FF4D781C1860407F49396109411C0C40367F7F084909496341490B18",
            INIT_RAM_17 => X"F0001F0F0018E00703000000FFF81FF8C0F81FF0FF0033300033008001F00000",
            INIT_RAM_18 => X"EE7A99E2972DB2E6B6ABD6224499B42B4A5BCE720CCBD5A114AFFFFFFAAAAAAB",
            INIT_RAM_19 => X"D318D9C482F8B719A5BECF0053B21095DB68C1F680194066381C4BB0CFFB3BED",
            INIT_RAM_1A => X"D8F5B2E70DDD89C19DC64440B486D3E5BBB4710805D45A72BEE2230CE1ED6C30",
            INIT_RAM_1B => X"6206211399B03840E27382229C3D6C4325FD24F6302666929D3DCC94B00A1CE7",
            INIT_RAM_1C => X"197AA1AEEC4FC1C825C7959C4C8ECBF66326933BABC8FDD46395B523A940D10F",
            INIT_RAM_1D => X"58AA836862292E136F55AD864D5B68B478988894F4B8E7AF44E146D54F4A2934",
            INIT_RAM_1E => X"772960E94C75A52717CDB34C133B32B126C3AC957C1D74AFEEEFAFFFBDFFCBEC",
            INIT_RAM_1F => X"AA973EC44266E64E8A1833A7AB5E234441F7F6E7266DF2AAE49D1F4DBF68934F",
            INIT_RAM_20 => X"1333FF40BFF2C1D9BD305E807EFA7F9540086F403FFD3DCAA0040B9413949B94",
            INIT_RAM_21 => X"C05A4AF64C174381002085A818210A0282888480316FF80787E66B6DBEDBEC57",
            INIT_RAM_22 => X"D17BA9EEA60083020C7005753054893445C8D8010D4CAD296622A44216125000",
            INIT_RAM_23 => X"75AF8FF5B681911A220C2F31AA11EF5F5B7FF7B5F0DB01E0835280ECDAD2F6EB",
            INIT_RAM_24 => X"4F104518D101DA011C1A0D0D1881428020228035A6B4D786EA27B6EB6DCBF7BB",
            INIT_RAM_25 => X"60C8620848E472C40C822490A7912194A1000630848E5881104340009110C4A1",
            INIT_RAM_26 => X"316034142EEA4292C29109702024158E7305DED75CC17660382860EDDDB10DDB",
            INIT_RAM_27 => X"002890C403B0908458100512A422416C0498924210883AFC892491009A249107",
            INIT_RAM_28 => X"A421299849E410F8F8C042A2100000A02608189080505114838924210B686287",
            INIT_RAM_29 => X"0600AEAC8C8D40939C322028781149BB9BBAA8D35C18B1085210472E8833391C",
            INIT_RAM_2A => X"F9C224CF927756663945235293239AD847CB89344AAD819AA29E5A6C7ADDCEA5",
            INIT_RAM_2B => X"84D22AB9D49CFEBCABA262CE0D408001A8091C110F55AE7BB9B1CE64D906C99C",
            INIT_RAM_2C => X"75BB65D96DADEB5D48B6B6B5AD8C559AE724C298CF3C6B690AC621378ACB0751",
            INIT_RAM_2D => X"9BDDB5D5A956B0DAD4338B04C38841AD106926663130EF0835A24D2666E9B5AD",
            INIT_RAM_2E => X"734C915B25B00C1F5D5C4C601648299D6720D7935D72465D99B26EBE4997666C",
            INIT_RAM_2F => X"C994C99708671280AE6AD43DD96DC940319CCE0904D76E7D976E7D926C508146",
            INIT_RAM_30 => X"4A12530688AA629E48D9CC81A88B6B2DAD09132224B211812E4F09E19A343542",
            INIT_RAM_31 => X"1327D55D6A20D6906530CB2201AB042C4F0B15A2B0C880231C0201A6100468C5",
            INIT_RAM_32 => X"7F7CF2C18354893901A629E71F51BFB6DB6B698601A1228185238A667B450A94",
            INIT_RAM_33 => X"00A9A10CC0133DAD24C5D99662AD2D4562CB6D5249365008C2A5AF56DDB198BE",
            INIT_RAM_34 => X"6A8126466D37E67D1430989CE0D80C2432835B0BC9A99882490492080950AACF",
            INIT_RAM_35 => X"0189014358935598F038B21A7957C4403B031243259091478A163104960908D2",
            INIT_RAM_36 => X"B12262CE66586B635306C4C6A64011B5885A2A4C41F381981ACCC0B5E1C124D2",
            INIT_RAM_37 => X"2ED0FCFA89B424F1A1859E665360062192435910DB4C210013404DA890035291",
            INIT_RAM_38 => X"146622A4690372F97223F3BBB8ABD18194141404141414141ECEE04F78EBDA3E",
            INIT_RAM_39 => X"0901030386D838BBCCE9DC01BEF18646552206B0D8A94ECC5C9034620C561810",
            INIT_RAM_3A => X"81D363427FC98CDC8D88233F5CCFE31222668F827196E0DC1B4B014A0E84386E",
            INIT_RAM_3B => X"984451C7FF36909224A112D8005093420494001000A65980DE253FFDA721BD99",
            INIT_RAM_3C => X"FFFFFFFFFFFEECFDADF95D273264DAB6E35B8AFE330021612525F2B410F9C9BF",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"A3FFB5B3792496DB65FF7FE693FB2CBEFFFFFFFFFFE7F3FF0000000000000000"
        )
        port map (
            DO => sdpb_inst_3_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_3_BLKSELA_i,
            BLKSELB => sdpb_inst_3_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_3_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_4: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"DA22DA1B031A8804A592014CD9ACD865020310241208912590482414B11104B4",
            INIT_RAM_01 => X"08478401030202400801180C2CCD00C06212016358E000008640050000080CEC",
            INIT_RAM_02 => X"C69D0A5008C2002904060000072E10244100058509A01026804114439504A08C",
            INIT_RAM_03 => X"4166049995828244D0A66D0862650B2C0010200206840320480145201120E340",
            INIT_RAM_04 => X"48422241A404057FC0C28CA995112A0CA502108249D0650A0CE542649589146C",
            INIT_RAM_05 => X"2422DC0423C8893024632031004012006904D2667229A3CA5010173491210082",
            INIT_RAM_06 => X"4A4AAA690220822AAA948809104CB0DA90151108826B4164600380091A360D24",
            INIT_RAM_07 => X"A42206360D0928033AEB688A8822B24194041036EC42104D0666A018404C24D0",
            INIT_RAM_08 => X"E13C202004670846222104C24A2207229114AB92084131408148A140A0404C40",
            INIT_RAM_09 => X"E006008349A22C6CA8C20420201942046246824810801081248C66165E4C2011",
            INIT_RAM_0A => X"0804D0082068180801248948248B0A0C80E304B6492C45A1254A592589112340",
            INIT_RAM_0B => X"11BB16704814068A040A400124A492D064110828888CD8014842338010A88251",
            INIT_RAM_0C => X"131810A228470404181A324915038200062340122264203B934024809258B103",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFF638DA25EFF5F74E11042284738C84E2245D4A20124933D22E",
            INIT_RAM_0E => X"04448B62B5ED800CB5A12514449998B08A631366D08D42096489024A8A091263",
            INIT_RAM_0F => X"FFB12124921442B319D684120A854F11248668EC16D86202281020559A340084",
            INIT_RAM_10 => X"7EFE415E7F59781C3060407F49192109410E06401C417F084109494141490B41",
            INIT_RAM_11 => X"51631436E42449497949451449517F49306008E03E1C633E044D186B14004F00",
            INIT_RAM_12 => X"0F78FFCCFF3E0073663CE0003F607E0303381CC00F07F000FF30060C18FF7E18",
            INIT_RAM_13 => X"0F0F1F00F0C0E00703000000FFF81FF8C0F81F00FF001FC000CC008001F0FF00",
            INIT_RAM_14 => X"7EFE415E7F74A0383060407F540424244404187F30807D04A47F544444445441",
            INIT_RAM_15 => X"51631436E42449497949451449517F49306008E03E1C633E044D186B14004F00",
            INIT_RAM_16 => X"3333FFCCFF59781C3060407F49192109410E06401C417F084109494141490B18",
            INIT_RAM_17 => X"0F0F1F00F030E00703000000FFF81FF8C0F81F00FF0066C000CC008001F0FF00",
            INIT_RAM_18 => X"0D44D1CC120D229400039400030D360280020428044201300280000003333330",
            INIT_RAM_19 => X"080084082081000011009B220830A22112102838344098020C6789264925A201",
            INIT_RAM_1A => X"9006C1B59C8C408428C24C042061C1B391882011182A8070B0C408C0E45CE984",
            INIT_RAM_1B => X"80630866466F16251063241461063231812601390101116CC18100119800C290",
            INIT_RAM_1C => X"3840CB11119B6430D99B2310040469B4C89A3044008E40005BA1302A37487200",
            INIT_RAM_1D => X"9918CB4CE46DA65A68419C31ED0442212330336361324D3580483322E84C0974",
            INIT_RAM_1E => X"219CE46DBC21B42000C000041519331000428061742C26BFEAEFEBFFB8EE31B0",
            INIT_RAM_1F => X"2010041830804220073909010F10C7002000E0133004D130604204001A60176D",
            INIT_RAM_20 => X"9777FF0ABFFD4CFBBB4F01A17EFD8461611940D2CF4AC272F2CEC14008C852C8",
            INIT_RAM_21 => X"853E1089961181092086D02D6C348B42828086102C04A537F7E983EFBED61397",
            INIT_RAM_22 => X"044E49392300020008606002D818331808136C01A10426894C02B01AD7121E50",
            INIT_RAM_23 => X"52961245149708A318004078C2214C29294290943666146113225B666A604A21",
            INIT_RAM_24 => X"4A035853650D28201490524024020490492492000008003000049390005A1083",
            INIT_RAM_25 => X"41424BC32954AAD54202492D246242739CE104BC32948AA8404D902485A54C14",
            INIT_RAM_26 => X"4215847EA2AA95521FD2A90BA5F415294D8729451361C3B0E243B09444999112",
            INIT_RAM_27 => X"61412D6A652939DC95683118A2A11A5549090421002B282DA2516BA51548EBA1",
            INIT_RAM_28 => X"A2108144B124928D0C375015A9B906230B9B352D5005530C3490421090129930",
            INIT_RAM_29 => X"736046622224A40809080A0017D7E922922AAB51562C5991518F40CD8005150A",
            INIT_RAM_2A => X"42B44D1424A0CCC9536865C52C442806B010509B92A0400B9690891002B36901",
            INIT_RAM_2B => X"0640069D1CE68D8040941400A12116D425B20122C054C4008C281149476B1231",
            INIT_RAM_2C => X"1DA5201315A5BB45C217B69DA294D44814C42992646122587634D32466281340",
            INIT_RAM_2D => X"20449954A3D2B256D8C429A198109C0C21148AC8986620939184229AC858BDA5",
            INIT_RAM_2E => X"6167485B6C9BA32020C1600AC4469920848E60944004C4C08804800018702201",
            INIT_RAM_2F => X"88446985678DE12290624421772204628B1804B259002A10302A113224C1880C",
            INIT_RAM_30 => X"849A5672E9B690940E2419954AA50CA08440844D8E448854C248330C21811984",
            INIT_RAM_31 => X"312575552AA80024881E644532A130C6483058066EB52AAB4B3199496B132D0A",
            INIT_RAM_32 => X"002B016BD7560452640941E5A031000000004342A415188408AC2E4000183B93",
            INIT_RAM_33 => X"CA42D20028002900CC99B167E54CA4C8A79FFC224921E800431CBC6366D00543",
            INIT_RAM_34 => X"19949230CCC5154279E63A60C8D1C46640812812C233150492492492A8020430",
            INIT_RAM_35 => X"4DB8FB23339008C2487B111B5AABEBBCD81524B065294ECBB0CC37E1CC12AF3B",
            INIT_RAM_36 => X"26B18CB601956E6608DCD330507ACCF145003E6CCD0B419630E8BCF1ECC71B73",
            INIT_RAM_37 => X"028101E0664108C4C6CFD51B681D8608890324C89A6375AB3346999F998E7302",
            INIT_RAM_38 => X"8199944A28745A00733222AAA8A04680C323332303030322116B200F73302423",
            INIT_RAM_39 => X"D692263A2AD9D9FAA36E0361BEE0608058DD547678750A720A64746C800198E7",
            INIT_RAM_3A => X"0614E5A8006323226795104254C822E0849A2074B60020040001AB03232D8291",
            INIT_RAM_3B => X"ECE4D144220251244925519B084011514AA114511609316963484008C9A2D0CC",
            INIT_RAM_3C => X"D369FFFFFFFEBC0786427448588978FB83640BB9921C2430DF277B12100141A1",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"F9B6C800068004929B2012136886D348FFFFFFFFFFF349FF0000000000000000"
        )
        port map (
            DO => sdpb_inst_4_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_4_BLKSELA_i,
            BLKSELB => sdpb_inst_4_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_4_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_5: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"9A0090D257E1E9F2020D35F80B580A89B87EA08040220482CE00804AD3B812E1",
            INIT_RAM_01 => X"6ADF3153685299DA432C6A794D9C90C8644A4D4B52E58065688C4A00D2AA8A88",
            INIT_RAM_02 => X"8C54D49B255F218DA558729229080912682EB2BDA360728D8108460487D542B9",
            INIT_RAM_03 => X"651C29A45622AA965AC71DB5DB15D34D2A86CAA6CC22944CD87B0C07B3D5873D",
            INIT_RAM_04 => X"2D6B3372B751416B0861D1365999DB51311B48CB6E1689A25176494D3750DA66",
            INIT_RAM_05 => X"ECAB13922352AD8569C6026256A5AB7EF2B5888C602AA08AF035B68CA535A6D1",
            INIT_RAM_06 => X"4C04B17E4936FBEFBCEEEEE598DD15ECE853376E66CD8EE77F510C02F06C1B01",
            INIT_RAM_07 => X"84BB8C2C1B3B1A3BEDB9E0DBEFBEFF7F273352A5CD739BBF3332CB45AD0D865F",
            INIT_RAM_08 => X"756EAA6A362FED6D9933C68453533FFFDDFFFB26CCF1A26CCFFFF5F13A3A3514",
            INIT_RAM_09 => X"92F14AA9667D98CA9DAE96CD91D8EA968FA459CD12DF9ADEA1B97D45675BD6E5",
            INIT_RAM_0A => X"08328A6DB7AD706D29B63D69B63D76B4C3D43CB6DB654584E5D97DB7DC97D36D",
            INIT_RAM_0B => X"BB11196064060C1364C909A086B4D3181494B414CD88895C695A604490A08041",
            INIT_RAM_0C => X"B7BF523BEAD9D859B0A3C4024DFF198168359754F9861B513960A49A8A26B4BD",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFFC6D9438808040410D7A91FCDA6E59AA2D4222E8C94B6692B6",
            INIT_RAM_0E => X"BF33725631A9BFF8E765614D8C9354AFB6C47ACDD3B24B2C8D9B7DA0A16B4913",
            INIT_RAM_0F => X"FFE324749A446AC6F9D4C640FAF46525555DDCC1B12499C0002ABFE54F9F523B",
            INIT_RAM_10 => X"3C0C417C7F710F777F3F7F016F7F3F7F7F7F7F7F7F60417F7F7F7F7F7F7F7E7F",
            INIT_RAM_11 => X"0341141C80006F7F037F67186373447F60000880083E411C007F332E7F070000",
            INIT_RAM_12 => X"077800CC181C004C7E7E00FF1F607E0303700EC01C003800FF30060C18005C18",
            INIT_RAM_13 => X"0F0F1800F0C0E0070300FF0018181800C018000000003FC000CC008001F0FF00",
            INIT_RAM_14 => X"3C0C417C7F64BC6C7C3C7C3F5C7C3CFC7C7C7C417FC0007FBC7E7C7C7C7F747F",
            INIT_RAM_15 => X"0341141C80006F7F037F67186373447F60000880083E411C007F332E7F070000",
            INIT_RAM_16 => X"993300CC18710F777F3F7F016F7F3F7F7F7F7F7F7F60417F7F7F7F7F7F7F7E18",
            INIT_RAM_17 => X"0F0F1800F078E0070300FF0018181800C01800000000CCC000CC008001F0FF00",
            INIT_RAM_18 => X"126D662BA7708653859085060EB6CB0A4202423A008A6AD80370000001696968",
            INIT_RAM_19 => X"A2B1218A297174F04A7CC1A8205888098DD08A0814020AC4824717A8193B8E2B",
            INIT_RAM_1A => X"65FC941EF7275B75926CCEC50DCC761EC6CADB457158C2122914631B15D636B1",
            INIT_RAM_1B => X"30C2090464E53C1576B5E146820C2C7207662CE11001132A6CD3DDA0EC4394CC",
            INIT_RAM_1C => X"AF458E511330310012002A500B19901E254C0BCC524B000111241D4BE2193A47",
            INIT_RAM_1D => X"2E2D35B3B832D3A5B462D744B28C48240060864E014125E760E842CD941D735B",
            INIT_RAM_1E => X"48E33136B6DADA6A35293499B64ECE254ABD090B83D74B1001000000462323D0",
            INIT_RAM_1F => X"E4643B08D49C4D89488C44C6CDA9818C138674A4D769CD40DB56D769A091B5B1",
            INIT_RAM_20 => X"0101F750C096FFF6F676848CC04800848484C24679BC02424242403FF3639363",
            INIT_RAM_21 => X"DE05736F043841B7DA55ACFAE86A7DB76F83ECC5E2A355700000336D96920000",
            INIT_RAM_22 => X"11CEBF3AFA183360CD9D16F4D0F14EB1B9DE086F53CE7C5EE20FC686BB7FBDE4",
            INIT_RAM_23 => X"738E46DD27F979B616C1007B9D35D43B0BC3B3B82CD682540E942056D7C5C663",
            INIT_RAM_24 => X"236B72C64BA718D057F75CFBB76A696D96D96D84708610D2740C93A9201E319E",
            INIT_RAM_25 => X"634FDC49BD5AAD5DCF7DD1B991B34A4A56B7DDC49BD69BB9EFB92ADB6E39E774",
            INIT_RAM_26 => X"4A5A9ADF44BD517D537E3EB3FC7E3BBDEB0F58C71CC3D661E8B4618CCC93A99B",
            INIT_RAM_27 => X"2C7D39CF35CD8D68E545ACAFFAADE31D493514631F5AAE4C2B45A2D9764F63D3",
            INIT_RAM_28 => X"431C3502A0ACFF48C9ABE3E73CE8B5952C8D3D3DD67D7967C75146319332DF3C",
            INIT_RAM_29 => X"C2EA059C2226DCF0F007070D2FFDFD2AD22FB85B64FDF3AAD30BE18AA046168B",
            INIT_RAM_2A => X"69B328C69030E5C6196120D19531980A43010BB74F6EA80CB447CF3B7F433D7F",
            INIT_RAM_2B => X"8021111C6355D44200010000121C08024204400C14D481718CD04820C384083C",
            INIT_RAM_2C => X"7D9FA523E48CFB15A836B23D8FE6F4F8C4ACBC9C790415753637A939DA79C3A1",
            INIT_RAM_2D => X"1D449AF18B5FD0D24504F83FA54A6BF1BE1487CF8FE9594D7E37C28FCF95B58C",
            INIT_RAM_2E => X"31C1218104154EA38673976794CBC9AEEC0A39E7F94CFCF98D687CAD1E7E634A",
            INIT_RAM_2F => X"997CF695E6DC9DFF67A1428CF763D8A888C56370B8FE6F4B3E6F5B3C4EBD51C6",
            INIT_RAM_30 => X"77FDAE2F944D50421563B8E3D330544B7FDBFC3D8E4311D6A5235F636D7E2EF4",
            INIT_RAM_31 => X"9E90AABAD4CDBFFD877664373308ABA5235EAF59114F6ECC6777BBBD6B6137BE",
            INIT_RAM_32 => X"DDD50640D2D3C466D468D67F668B4DB6DB6F5134F5DF2F91DFDD59BDBFEFC476",
            INIT_RAM_33 => X"200000400003A52382B0344174F7FE29030DB8C00017A00003939FE76E988F55",
            INIT_RAM_34 => X"B5F6DB927AE19562B1CF7E4459F5852D2D530AD88A60A4349B2936541356A000",
            INIT_RAM_35 => X"E7DED197FFF370BB653614BEFEEABAB819001266288C6CA1616F6AC07F40FE7E",
            INIT_RAM_36 => X"1D6B0865E40FF7DFD9FFF6439A5F2E7CC84A46DFF8C02BC53C3E1A7872EFF236",
            INIT_RAM_37 => X"22D441F0B21CC7D158ADB412A62E2D70A71E8EA5BEDCFF7EFFF24F5BB6D7BD7E",
            INIT_RAM_38 => X"F39F928197A3A2FF84CDD444431F8005A141414141010160125E596A5E240555",
            INIT_RAM_39 => X"CC78F8FF21B515B682578B8B6DB8D21083B75D7F3DE79E54C7413CD87221E2F7",
            INIT_RAM_3A => X"7CE6773C8681657777D5352AC7E03E2816322762AC94BE97D2D37EBFC64CC464",
            INIT_RAM_3B => X"4AEE71C7E0A3349300567DF5E59CE2F3CFA77DFDDEEDB17D46BD043E8D7A9FBA",
            INIT_RAM_3C => X"D349FFFFFFFEE6FCC403CD4A5ECDC99E05499A78B6206049842CF6247BF8E8DF",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"FDA249B6948DB249926DB4986D2492407FFFFFFFFFF209FF0000000000000000"
        )
        port map (
            DO => sdpb_inst_5_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_5_BLKSELA_i,
            BLKSELB => sdpb_inst_5_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_5_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_6: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"0AAA4900011644062659432A908A90031101022512888124304A253118004191",
            INIT_RAM_01 => X"423791D44410B42128C52A5D0406245228A09408020A250C2021984A081A6000",
            INIT_RAM_02 => X"A500C42018555C2050C31000242805910000084D012F3004803048121344480A",
            INIT_RAM_03 => X"510EE00A14600885510E8D10928540008544EBA2A42880100053AE1308A0A298",
            INIT_RAM_04 => X"385AAA88A910056AA0C2C02411555B0061FA36A36ADE0303000446000480915D",
            INIT_RAM_05 => X"A42428646C108A2D08F70068081A04806066E21C620A8182D00610D523E279BE",
            INIT_RAM_06 => X"4C4C1220109841041188008B44738D2211A00018031499196A78D02010242900",
            INIT_RAM_07 => X"D60084240929284B45131E610410448BC040116800C0064116D844121050A8A2",
            INIT_RAM_08 => X"C598B230593248874CC200D8C008204400484780208060020891001A05454772",
            INIT_RAM_09 => X"4D2C30C293334E7C88C4687242444068331524701124E12478D4762E6CEC24B6",
            INIT_RAM_0A => X"401697CB2C2BBBC00125635525635458AAC3EFDB6DB6DF237962712509698A92",
            INIT_RAM_0B => X"55D5D6AF4BD404E0040A4B1F74A492D7C48643E3BAEFAF2548523A0204081210",
            INIT_RAM_0C => X"1A1210AC28434D0E9A0B509005404AC083832914CCF4403F554024B175C88641",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFFD299B868281434318544E2C560D4FF2F63DDF0174F1A39763",
            INIT_RAM_0E => X"2155764CB5A91FF8A52121043C9332A28A430624B0A946D0B489368282C90940",
            INIT_RAM_0F => X"FFE1B7C5F20640925095841A20B84299450CE93E46DB661F3FB02065FAB40062",
            INIT_RAM_10 => X"18080068006107637F1F3F01267F1E7F3E7F7F7F7F20007F3E7F7F7F3E7F7C3E",
            INIT_RAM_11 => X"0241140800002636033E27182262403E40000800082A0000003263247F070000",
            INIT_RAM_12 => X"031000331808000C3CE700FF0E603C03FFE007FF180018000030060C18001818",
            INIT_RAM_13 => X"0F0F1800F0C0E0070300FFFF18181800C018000000007F300033FF8001F0FF00",
            INIT_RAM_14 => X"1808006800449C441C1C3C04487C18FC387C7C007F40007F98083838387F203E",
            INIT_RAM_15 => X"0241140800002636033E27182262403E40000800082A0000003263247F070000",
            INIT_RAM_16 => X"CCCC0033186107637F1F3F01267F1E7F3E7F7F7F7F20007F3E7F7F7F3E7F7C18",
            INIT_RAM_17 => X"0F0F1800F078E0070300FFFF18181800C0180000000099300033FF8001F0FF00",
            INIT_RAM_18 => X"321A9ABF8115B49582AA52A54ABD2640109014AA100035355100000005B24DB0",
            INIT_RAM_19 => X"C398D16C355D954996969E19C3A4B014527C1D5E875C64A2292BC4A2E92BAA2D",
            INIT_RAM_1A => X"997EF1F5A9D91A990C8B66B2F54C95F53B2EA2CCB5C501489742421D65084821",
            INIT_RAM_1B => X"242D6AD5557C5285AA94659409446284AB24775CF849469FDDB95415DA91DC22",
            INIT_RAM_1C => X"9313AD377556E5ACBD57B6C54496CFE0C622AA55ADAEAC0153112D01ABC83A9E",
            INIT_RAM_1D => X"FBFED24C6379AC9A4B55898669C502816AAC2AF6F9B8CF652942127F6BCB5624",
            INIT_RAM_1E => X"65AD45ED68A7B5CB2588A554E19337A04860A9142E0C26BBBFAAAAAABB980EAE",
            INIT_RAM_1F => X"6AA72CE6862E8A0EEB116B253A77B2480B75C0B5B54978BAB59554281F69626F",
            INIT_RAM_20 => X"0101F70026600000000000A033337F7B7B3B00500001BDBDBD9DA13BB2958094",
            INIT_RAM_21 => X"8C4C39A3C695A1124CE1304B4D2C12DBB48134AC4115EED000038F6D96920000",
            INIT_RAM_22 => X"A4CE1B386B48122048A64B279A30365EDC538D316A07C71B0C04C6541F26D0C4",
            INIT_RAM_23 => X"1086524801A1B00FE040FF86F8219C2909C29299B6433DE3F303DF6241714261",
            INIT_RAM_24 => X"48235A437945086003AE0FD711200BA6BA6BA6A1142A85649824938249061284",
            INIT_RAM_25 => X"06C4F1411168B4004134B4902428008421026F141114A008269DE469A5BDAB37",
            INIT_RAM_26 => X"002D2A5D2C15013503303A8A604C6B38C9A708410269C934E61B3494CC998440",
            INIT_RAM_27 => X"711805AD5174A0023D8A0506D6E0C044401124842D1204C82050024CA7250246",
            INIT_RAM_28 => X"0847381822C6747071024196B54540A04552848058F5D9058112484281EA0A95",
            INIT_RAM_29 => X"6F01F606AAED6C1A156666446BB5D80000015708267CF98001BEC8A200725A2D",
            INIT_RAM_2A => X"0A956910A4A4CAA953A874C52C552890855210911645C22AF290B94D3E7BE9ED",
            INIT_RAM_2B => X"52FAA4F5494E9819F7FCFDFDEDE3F7FDBDF3BFE3EAD4A82B2953944D930953A1",
            INIT_RAM_2C => X"56D141697EC6ADAE929ADB16C0B8C79E41241042CF3D4D3241C1B088CBEF1679",
            INIT_RAM_2D => X"93EEDA9AC16C1267E85503F9E19C01101145AEEEBE784F00320228AEEEF0D6C6",
            INIT_RAM_2E => X"00E4808000015628081F392400410461B4B6E5A73C5E5E5C891E4E2F5AB72A57",
            INIT_RAM_2F => X"083452806CEE913110A2C421BF6365A0A80100789DC72256B72A469408304080",
            INIT_RAM_30 => X"44D487244544169084589DC140044B090C42C54FA6D40085DE4813E1A0201910",
            INIT_RAM_31 => X"3B24088C6000C424A856ED42000F25DE48130980400D0004210080CA10356BD6",
            INIT_RAM_32 => X"FDDFDE0000028F1B6482496B8F21A0000005639064090684084FA0A6A2013762",
            INIT_RAM_33 => X"DF7EFFBFFC03A100A31541758044848BD7D7B0700003E80801FB936B6E9005F7",
            INIT_RAM_34 => X"11D7FF304C757300D5E6F2EC68909C4458810992122A951000200044020407BD",
            INIT_RAM_35 => X"6F9CF042108033C0D01A721B12AAAFFCE6FFA4B741294585A644314D5412AADA",
            INIT_RAM_36 => X"AC30EEAE03D54A621BC496CD162E5DE100000A4CEDEB811692A89D65458536D2",
            INIT_RAM_37 => X"0A013C88292C60F56FCCD05A134CA43393431DD09A60B52F3A660982908212C3",
            INIT_RAM_38 => X"81FC83F9790522016110800080A01180AA8A8A8A8AAAAA8AB7E7000C47719501",
            INIT_RAM_39 => X"9632651BACD9F99A0B60D329A6C1648413B15436B0F7C48ED6D5646A05DD801F",
            INIT_RAM_3A => X"85E5C7E8029898AAEB151D019488251E74B6AF74B580200400052F620B099CB8",
            INIT_RAM_3B => X"7C82A083D586940100445898A08882334E2334C91649A839731513E9E9A2E098",
            INIT_RAM_3C => X"B7FFFFFFFFFEF5AEAEABE54A50A96BC3076E8B34A3F225408F0662A031A8A05E",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"BB2DBC936DE49249B6FB6FB6DB7DFFDEFFFFFFFFFFFFF7FF0000000000000000"
        )
        port map (
            DO => sdpb_inst_6_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_6_BLKSELA_i,
            BLKSELB => sdpb_inst_6_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_6_DI_i,
            ADB => adb(13 downto 0)
        );

    sdpb_inst_7: SDPB
        generic map (
            READ_MODE => '0',
            BIT_WIDTH_0 => 1,
            BIT_WIDTH_1 => 1,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"DAAAD91B573ECC56B51DE66ADBBADAEF2B167F379BCC89B6B26F37B3A3BB97B5",
            INIT_RAM_01 => X"5B67ED1E7896E4736BCD6A6F699F369B4CF0D96B5ACF37294EE4526318BAECEC",
            INIT_RAM_02 => X"49155EE37B58E1AD621A6C4905E202D1E04E3CE16550C19543E63982F594184A",
            INIT_RAM_03 => X"19E6EDAB911A4AE543B6EC2532E41B6DCC567234C8D2D770DF894410B315D685",
            INIT_RAM_04 => X"1903A8DA8C14406FBB019DBD11DC1B5DE57B76F360D6EF2A5DE66E6DB73F8655",
            INIT_RAM_05 => X"AD2C8AE7BD5CA239EE7FFBAB5CB32CCAE2C4DBC56BAA9DAAA0572AF2BA676D36",
            INIT_RAM_06 => X"69214704A445145145A955562ABBAB85668AAAB95552322A5C23BBC4B42D2B42",
            INIT_RAM_07 => X"AD556D2D0B6B6B929052395555554EABD4AAAB2AA5C94C82A5DD0E5739752AEC",
            INIT_RAM_08 => X"E79CF373A873258B46EE75DA0A4AA9552AAB57D2AB9D694AAAD54AA8A5555555",
            INIT_RAM_09 => X"5D35F6DA91774CFCA5CD68F34C952968B36534D14BA7A3A3B1CD76664E6CC6F6",
            INIT_RAM_0A => X"00024CC71CE65FC9D492E73892E7353871CFE6DB6DB7FF9630E1589394A3B293",
            INIT_RAM_0B => X"555D43FC0B11CE6A52A5263A607208CC5257674CAAAAEAF105297974C2040908",
            INIT_RAM_0C => X"3B394A9E562ABD3E7A7B3B6D9C176AFBDAA7CC4EEED19277F71C9263248A5765",
            INIT_RAM_0D => X"FFFFFFFFFFFFFFF354B8EC02010302DEA8B012BDAA92F2B6000216A463975777",
            INIT_RAM_0E => X"BB77D6CEB5A9BFEAED69694775B5F4AEBAD49EA5D7C86BD81CA974C3A2894043",
            INIT_RAM_0F => X"FFAFFF67B346C89295A4B553D894473175D4E160A0000010400FDF99F1E3FABB",
            INIT_RAM_10 => X"0000004000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_11 => X"0000000000000000000000000000000000000000000800000000000014000000",
            INIT_RAM_12 => X"010000331800000000C3000000600003FFC003FF180018000030060C18000018",
            INIT_RAM_13 => X"0F0F1800F0C0E0070300FFFF18181800C01800000000FF300033FF8001F0FF00",
            INIT_RAM_14 => X"0000004000000000000000040000000000000000000000000000000000000000",
            INIT_RAM_15 => X"0000000000000000000000000000000000000000000800000000000014000000",
            INIT_RAM_16 => X"66CC003318000000000000000000000000000000000000000000000000000018",
            INIT_RAM_17 => X"0F0F1800F000E0070300FFFF18181800C0180000000033300033FF8001F0FF00",
            INIT_RAM_18 => X"672FD07F93209252C3FEF7F7EFBDB4294E494E5FCEE95FA7FA500000063C71C0",
            INIT_RAM_19 => X"EB8DC16F3829E79CD4EBDF13E9F03B1473669EB3D74EE6F71DEFCDCBEB7D8EA7",
            INIT_RAM_1A => X"D1F7F5E3B9995BC9288F6EF2E5ED9737332EF3DCDDFFE1DFBB67625E4118EC25",
            INIT_RAM_1B => X"72A5295555500255FFBDB5D6A92D2A42A56D1B1D6C21572F8703FEB1F34ADE77",
            INIT_RAM_1C => X"3838AD55555745AEBF973A8FECDCE9B0CAA62B75F6FF57FE38149729EB5DBBC6",
            INIT_RAM_1D => X"FBFFD34CE77DB69A6DFF99D6E9AD2A9D72EEAEFAE1F2AA2D4420D2FFEDCF6464",
            INIT_RAM_1E => X"B3BDC5EDB8F7B68DB6CF379E4513A3B56EC5CDBE345974BAAFFAFEABA8AB2A36",
            INIT_RAM_1F => X"BFC7B66ED673AE2F3F316B37BE7BB66C0486B2F5246D51E2A6DF9E4F3A4DC66D",
            INIT_RAM_20 => X"0311F7DB634EF6FFFF7FFFE921A77B7B7B3B7FC00042000000001E3E9BDEC1DE",
            INIT_RAM_21 => X"99A4764DD6ABE9334CE676EF6D7C59D9B623B35684000007FCC80B6F97B21010",
            INIT_RAM_22 => X"155E3978E3522648991C275F9AD17E3DD99F8D73676B6F7A2A8E1B185236C299",
            INIT_RAM_23 => X"75BA9251B7338DD3FA910000F965052B4A52B6A0365700600320006250F656AA",
            INIT_RAM_24 => X"4F73FF57F9A55AC45D34579A3673792492492435E6BCD6B6D88DB78B6D92B5B9",
            INIT_RAM_25 => X"726E9969B9DEEF7FFBA499BDA7BB6BFFFFF769969B9EDFFF748FE6C937BDEF9C",
            INIT_RAM_26 => X"6B5C225788E18071827018C0E01D0318C9AF1AD75A6BC535E23B35AD55B9899B",
            INIT_RAM_27 => X"7D79BDEF77ED9CEAF76F952E9BBDC27FEDB1B6F7B9A3B881235180EDC76E00E4",
            INIT_RAM_28 => X"CF7ED0F6EBEC2666E693FBB7BDFDF2A46DCB95B176B773E5851B6F7BDBB2CF1C",
            INIT_RAM_29 => X"EF68062EAAAEE77A716E6E6C4AF579B3DB3EABF3CE7CF98AFBBBCDAEA04477BB",
            INIT_RAM_2A => X"9B166DD9B6F6EAAD7BAD76D734673AD8859B12951B0CCBBFB29EFD5C7B7AC5ED",
            INIT_RAM_2B => X"F2CFF7C46E4E14A2040101010000002000044008007DAD62390C18491B895B39",
            INIT_RAM_2C => X"77E9BDA177EFEFD78A9EFFB7FCE65E8C93CEB1CAEC61703177B2F3917F6D174D",
            INIT_RAM_2D => X"3B7FFC7DE9731A777555DDEF2B186527B155CE8EDBCAC90CB4F62AAE8ED0F7EF",
            INIT_RAM_2E => X"3964FD09249DFA29AE5B2E4CD2EB1CA6A0AABB875B6C4C5BEDA8EDBD0A16F36A",
            INIT_RAM_2F => X"5D66F0D3EEE8B1E3132AD4BD276BC522A9CE67E2F1DEFB6A16F36A1378F1DD67",
            INIT_RAM_30 => X"C79C7C64ADF4569ED7E7D9DDEFF7E4FD3DCD9E7DAEE7DC7CFE4F5E072CA7BF62",
            INIT_RAM_31 => X"3B27BFEDEFFD9CE4CFAEEE71BBFCBAFE4F5F2F93DA7DBFFBD777BAF9FF757FDE",
            INIT_RAM_32 => X"5D5552E9D2FBE41344E24DB1831389249249E2E4E4DDACD4D8C99324AE653FC6",
            INIT_RAM_33 => X"00000000000335A7A6B5F4F3D2C6D2EBF5D7FEF249340808019BB777FFBAAF57",
            INIT_RAM_34 => X"39DC923AE8C39DEAD5AEF3ECED91DC2C317B4B19FB6934A24944928BBDFBF000",
            INIT_RAM_35 => X"6F9CF96639DE5BCA991B733B32AAAFAE000012762C9CEEC9B7EE63ECFE49FF73",
            INIT_RAM_36 => X"9CF3AA76F74FCF477BEE9F6FD65F5D66EFFF7F6DECE9CB0EBA7C5D64C58FBB7B",
            INIT_RAM_37 => X"87DD01B42A55A7D467CFDD1E3B2EAC5B9B831ED99A67E7BE7A475D1FDBDF7A8E",
            INIT_RAM_38 => X"773156260C88D0788401459D10006E19020216060302020213E3A97FFBF8277B",
            INIT_RAM_39 => X"0AF9F7DE2791F1F3A3C5CBAB3CFCE252FB6BFE66B1F8144ECEE562CC861E00A0",
            INIT_RAM_3A => X"7E07C7E882AAAAAAEB1FB84106843152A67B2452E6D2664CC94BBE4667EDF85C",
            INIT_RAM_3B => X"FCEEF9E7EA2B9892249FF1D16F16FB9BEF35FFE7FE8DA97DE7605018CFA3C989",
            INIT_RAM_3C => X"DA4DFFFFFFFEBE57E7527E6C78CDFCFF81FF4FEAB417357DADAFDEB75A51C99F",
            INIT_RAM_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_RAM_3F => X"FD64980126800000926926D24924DA497FFFFFFFFFF34DFF0000000000000000"
        )
        port map (
            DO => sdpb_inst_7_DO_o,
            CLKA => clka,
            CEA => cea,
            CLKB => clkb,
            CEB => ceb,
            OCE => oce,
            RESET => reset,
            BLKSELA => sdpb_inst_7_BLKSELA_i,
            BLKSELB => sdpb_inst_7_BLKSELB_i,
            ADA => ada(13 downto 0),
            DI => sdpb_inst_7_DI_i,
            ADB => adb(13 downto 0)
        );

end Behavioral; --Gowin_SDPB_kernal_rom_16k_gw5a
